# original pdn
.title 20200622-104926
.option rshunt = 1.0e12
.subckt PcbBuckConverter VDD VSS
C1 VDD 12 2340uF
R1 12 13 0Ohm
L1 13 VSS 0nH
C2 VDD 22 0uF
R2 22 23 1000000000000.0Ohm
L2 23 VSS 0nH
Ls VDD 31 0.33uH
Rs 31 32 20mOhm
Vs 32 VSS 1.1
.ends PcbBuckConverter

.subckt PcbModelLumped VDD1 VSS1 VDD2 VSS2
Rs1 VDD1 11 1000mOhm
Ls1 11 VDD2 0nH
Rs2 VSS1 21 1000mOhm
Ls2 21 VSS2 0nH
Rp VDD2 VDD2M 0mOhm
Cp VDD2M VSS2 0uF
.ends PcbModelLumped

.subckt dut VDD VSS
R_X10Y10VDD_X20Y10VDD X10Y10VDD X15Y10VDD 25mOhm
L_X10Y10VDD_X20Y10VDD X15Y10VDD X20Y10VDD 2.91e-06nH
R_X10Y10VSS_X20Y10VSS X10Y10VSS X15Y10VSS 25mOhm
L_X10Y10VSS_X20Y10VSS X15Y10VSS X20Y10VSS 2.91e-06nH
R_X20Y10VDD_X30Y10VDD X20Y10VDD X25Y10VDD 25mOhm
L_X20Y10VDD_X30Y10VDD X25Y10VDD X30Y10VDD 2.91e-06nH
R_X20Y10VSS_X30Y10VSS X20Y10VSS X25Y10VSS 25mOhm
L_X20Y10VSS_X30Y10VSS X25Y10VSS X30Y10VSS 2.91e-06nH
R_X30Y10VDD_X40Y10VDD X30Y10VDD X35Y10VDD 25mOhm
L_X30Y10VDD_X40Y10VDD X35Y10VDD X40Y10VDD 2.91e-06nH
R_X30Y10VSS_X40Y10VSS X30Y10VSS X35Y10VSS 25mOhm
L_X30Y10VSS_X40Y10VSS X35Y10VSS X40Y10VSS 2.91e-06nH
R_X40Y10VDD_X50Y10VDD X40Y10VDD X45Y10VDD 25mOhm
L_X40Y10VDD_X50Y10VDD X45Y10VDD X50Y10VDD 2.91e-06nH
R_X40Y10VSS_X50Y10VSS X40Y10VSS X45Y10VSS 25mOhm
L_X40Y10VSS_X50Y10VSS X45Y10VSS X50Y10VSS 2.91e-06nH
R_X50Y10VDD_X60Y10VDD X50Y10VDD X55Y10VDD 25mOhm
L_X50Y10VDD_X60Y10VDD X55Y10VDD X60Y10VDD 2.91e-06nH
R_X50Y10VSS_X60Y10VSS X50Y10VSS X55Y10VSS 25mOhm
L_X50Y10VSS_X60Y10VSS X55Y10VSS X60Y10VSS 2.91e-06nH
R_X60Y10VDD_X70Y10VDD X60Y10VDD X65Y10VDD 25mOhm
L_X60Y10VDD_X70Y10VDD X65Y10VDD X70Y10VDD 2.91e-06nH
R_X60Y10VSS_X70Y10VSS X60Y10VSS X65Y10VSS 25mOhm
L_X60Y10VSS_X70Y10VSS X65Y10VSS X70Y10VSS 2.91e-06nH
R_X70Y10VDD_X80Y10VDD X70Y10VDD X75Y10VDD 25mOhm
L_X70Y10VDD_X80Y10VDD X75Y10VDD X80Y10VDD 2.91e-06nH
R_X70Y10VSS_X80Y10VSS X70Y10VSS X75Y10VSS 25mOhm
L_X70Y10VSS_X80Y10VSS X75Y10VSS X80Y10VSS 2.91e-06nH
R_X80Y10VDD_X90Y10VDD X80Y10VDD X85Y10VDD 25mOhm
L_X80Y10VDD_X90Y10VDD X85Y10VDD X90Y10VDD 2.91e-06nH
R_X80Y10VSS_X90Y10VSS X80Y10VSS X85Y10VSS 25mOhm
L_X80Y10VSS_X90Y10VSS X85Y10VSS X90Y10VSS 2.91e-06nH
R_X90Y10VDD_X100Y10VDD X90Y10VDD X95Y10VDD 25mOhm
L_X90Y10VDD_X100Y10VDD X95Y10VDD X100Y10VDD 2.91e-06nH
R_X90Y10VSS_X100Y10VSS X90Y10VSS X95Y10VSS 25mOhm
L_X90Y10VSS_X100Y10VSS X95Y10VSS X100Y10VSS 2.91e-06nH
R_X100Y10VDD_X110Y10VDD X100Y10VDD X105Y10VDD 25mOhm
L_X100Y10VDD_X110Y10VDD X105Y10VDD X110Y10VDD 2.91e-06nH
R_X100Y10VSS_X110Y10VSS X100Y10VSS X105Y10VSS 25mOhm
L_X100Y10VSS_X110Y10VSS X105Y10VSS X110Y10VSS 2.91e-06nH
R_X110Y10VDD_X120Y10VDD X110Y10VDD X115Y10VDD 25mOhm
L_X110Y10VDD_X120Y10VDD X115Y10VDD X120Y10VDD 2.91e-06nH
R_X110Y10VSS_X120Y10VSS X110Y10VSS X115Y10VSS 25mOhm
L_X110Y10VSS_X120Y10VSS X115Y10VSS X120Y10VSS 2.91e-06nH
R_X10Y20VDD_X20Y20VDD X10Y20VDD X15Y20VDD 25mOhm
L_X10Y20VDD_X20Y20VDD X15Y20VDD X20Y20VDD 2.91e-06nH
R_X10Y20VSS_X20Y20VSS X10Y20VSS X15Y20VSS 25mOhm
L_X10Y20VSS_X20Y20VSS X15Y20VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X30Y20VDD X20Y20VDD X25Y20VDD 25mOhm
L_X20Y20VDD_X30Y20VDD X25Y20VDD X30Y20VDD 2.91e-06nH
R_X20Y20VSS_X30Y20VSS X20Y20VSS X25Y20VSS 25mOhm
L_X20Y20VSS_X30Y20VSS X25Y20VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X40Y20VDD X30Y20VDD X35Y20VDD 25mOhm
L_X30Y20VDD_X40Y20VDD X35Y20VDD X40Y20VDD 2.91e-06nH
R_X30Y20VSS_X40Y20VSS X30Y20VSS X35Y20VSS 25mOhm
L_X30Y20VSS_X40Y20VSS X35Y20VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X50Y20VDD X40Y20VDD X45Y20VDD 25mOhm
L_X40Y20VDD_X50Y20VDD X45Y20VDD X50Y20VDD 2.91e-06nH
R_X40Y20VSS_X50Y20VSS X40Y20VSS X45Y20VSS 25mOhm
L_X40Y20VSS_X50Y20VSS X45Y20VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X60Y20VDD X50Y20VDD X55Y20VDD 25mOhm
L_X50Y20VDD_X60Y20VDD X55Y20VDD X60Y20VDD 2.91e-06nH
R_X50Y20VSS_X60Y20VSS X50Y20VSS X55Y20VSS 25mOhm
L_X50Y20VSS_X60Y20VSS X55Y20VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X70Y20VDD X60Y20VDD X65Y20VDD 25mOhm
L_X60Y20VDD_X70Y20VDD X65Y20VDD X70Y20VDD 2.91e-06nH
R_X60Y20VSS_X70Y20VSS X60Y20VSS X65Y20VSS 25mOhm
L_X60Y20VSS_X70Y20VSS X65Y20VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X80Y20VDD X70Y20VDD X75Y20VDD 25mOhm
L_X70Y20VDD_X80Y20VDD X75Y20VDD X80Y20VDD 2.91e-06nH
R_X70Y20VSS_X80Y20VSS X70Y20VSS X75Y20VSS 25mOhm
L_X70Y20VSS_X80Y20VSS X75Y20VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X90Y20VDD X80Y20VDD X85Y20VDD 25mOhm
L_X80Y20VDD_X90Y20VDD X85Y20VDD X90Y20VDD 2.91e-06nH
R_X80Y20VSS_X90Y20VSS X80Y20VSS X85Y20VSS 25mOhm
L_X80Y20VSS_X90Y20VSS X85Y20VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X100Y20VDD X90Y20VDD X95Y20VDD 25mOhm
L_X90Y20VDD_X100Y20VDD X95Y20VDD X100Y20VDD 2.91e-06nH
R_X90Y20VSS_X100Y20VSS X90Y20VSS X95Y20VSS 25mOhm
L_X90Y20VSS_X100Y20VSS X95Y20VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X110Y20VDD X100Y20VDD X105Y20VDD 25mOhm
L_X100Y20VDD_X110Y20VDD X105Y20VDD X110Y20VDD 2.91e-06nH
R_X100Y20VSS_X110Y20VSS X100Y20VSS X105Y20VSS 25mOhm
L_X100Y20VSS_X110Y20VSS X105Y20VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X120Y20VDD X110Y20VDD X115Y20VDD 25mOhm
L_X110Y20VDD_X120Y20VDD X115Y20VDD X120Y20VDD 2.91e-06nH
R_X110Y20VSS_X120Y20VSS X110Y20VSS X115Y20VSS 25mOhm
L_X110Y20VSS_X120Y20VSS X115Y20VSS X120Y20VSS 2.91e-06nH
R_X10Y30VDD_X20Y30VDD X10Y30VDD X15Y30VDD 25mOhm
L_X10Y30VDD_X20Y30VDD X15Y30VDD X20Y30VDD 2.91e-06nH
R_X10Y30VSS_X20Y30VSS X10Y30VSS X15Y30VSS 25mOhm
L_X10Y30VSS_X20Y30VSS X15Y30VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X30Y30VDD X20Y30VDD X25Y30VDD 25mOhm
L_X20Y30VDD_X30Y30VDD X25Y30VDD X30Y30VDD 2.91e-06nH
R_X20Y30VSS_X30Y30VSS X20Y30VSS X25Y30VSS 25mOhm
L_X20Y30VSS_X30Y30VSS X25Y30VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X40Y30VDD X30Y30VDD X35Y30VDD 25mOhm
L_X30Y30VDD_X40Y30VDD X35Y30VDD X40Y30VDD 2.91e-06nH
R_X30Y30VSS_X40Y30VSS X30Y30VSS X35Y30VSS 25mOhm
L_X30Y30VSS_X40Y30VSS X35Y30VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X50Y30VDD X40Y30VDD X45Y30VDD 25mOhm
L_X40Y30VDD_X50Y30VDD X45Y30VDD X50Y30VDD 2.91e-06nH
R_X40Y30VSS_X50Y30VSS X40Y30VSS X45Y30VSS 25mOhm
L_X40Y30VSS_X50Y30VSS X45Y30VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X60Y30VDD X50Y30VDD X55Y30VDD 25mOhm
L_X50Y30VDD_X60Y30VDD X55Y30VDD X60Y30VDD 2.91e-06nH
R_X50Y30VSS_X60Y30VSS X50Y30VSS X55Y30VSS 25mOhm
L_X50Y30VSS_X60Y30VSS X55Y30VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X70Y30VDD X60Y30VDD X65Y30VDD 25mOhm
L_X60Y30VDD_X70Y30VDD X65Y30VDD X70Y30VDD 2.91e-06nH
R_X60Y30VSS_X70Y30VSS X60Y30VSS X65Y30VSS 25mOhm
L_X60Y30VSS_X70Y30VSS X65Y30VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X80Y30VDD X70Y30VDD X75Y30VDD 25mOhm
L_X70Y30VDD_X80Y30VDD X75Y30VDD X80Y30VDD 2.91e-06nH
R_X70Y30VSS_X80Y30VSS X70Y30VSS X75Y30VSS 25mOhm
L_X70Y30VSS_X80Y30VSS X75Y30VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X90Y30VDD X80Y30VDD X85Y30VDD 25mOhm
L_X80Y30VDD_X90Y30VDD X85Y30VDD X90Y30VDD 2.91e-06nH
R_X80Y30VSS_X90Y30VSS X80Y30VSS X85Y30VSS 25mOhm
L_X80Y30VSS_X90Y30VSS X85Y30VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X100Y30VDD X90Y30VDD X95Y30VDD 25mOhm
L_X90Y30VDD_X100Y30VDD X95Y30VDD X100Y30VDD 2.91e-06nH
R_X90Y30VSS_X100Y30VSS X90Y30VSS X95Y30VSS 25mOhm
L_X90Y30VSS_X100Y30VSS X95Y30VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X110Y30VDD X100Y30VDD X105Y30VDD 25mOhm
L_X100Y30VDD_X110Y30VDD X105Y30VDD X110Y30VDD 2.91e-06nH
R_X100Y30VSS_X110Y30VSS X100Y30VSS X105Y30VSS 25mOhm
L_X100Y30VSS_X110Y30VSS X105Y30VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X120Y30VDD X110Y30VDD X115Y30VDD 25mOhm
L_X110Y30VDD_X120Y30VDD X115Y30VDD X120Y30VDD 2.91e-06nH
R_X110Y30VSS_X120Y30VSS X110Y30VSS X115Y30VSS 25mOhm
L_X110Y30VSS_X120Y30VSS X115Y30VSS X120Y30VSS 2.91e-06nH
R_X10Y40VDD_X20Y40VDD X10Y40VDD X15Y40VDD 25mOhm
L_X10Y40VDD_X20Y40VDD X15Y40VDD X20Y40VDD 2.91e-06nH
R_X10Y40VSS_X20Y40VSS X10Y40VSS X15Y40VSS 25mOhm
L_X10Y40VSS_X20Y40VSS X15Y40VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X30Y40VDD X20Y40VDD X25Y40VDD 25mOhm
L_X20Y40VDD_X30Y40VDD X25Y40VDD X30Y40VDD 2.91e-06nH
R_X20Y40VSS_X30Y40VSS X20Y40VSS X25Y40VSS 25mOhm
L_X20Y40VSS_X30Y40VSS X25Y40VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X40Y40VDD X30Y40VDD X35Y40VDD 25mOhm
L_X30Y40VDD_X40Y40VDD X35Y40VDD X40Y40VDD 2.91e-06nH
R_X30Y40VSS_X40Y40VSS X30Y40VSS X35Y40VSS 25mOhm
L_X30Y40VSS_X40Y40VSS X35Y40VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X50Y40VDD X40Y40VDD X45Y40VDD 25mOhm
L_X40Y40VDD_X50Y40VDD X45Y40VDD X50Y40VDD 2.91e-06nH
R_X40Y40VSS_X50Y40VSS X40Y40VSS X45Y40VSS 25mOhm
L_X40Y40VSS_X50Y40VSS X45Y40VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X60Y40VDD X50Y40VDD X55Y40VDD 25mOhm
L_X50Y40VDD_X60Y40VDD X55Y40VDD X60Y40VDD 2.91e-06nH
R_X50Y40VSS_X60Y40VSS X50Y40VSS X55Y40VSS 25mOhm
L_X50Y40VSS_X60Y40VSS X55Y40VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X70Y40VDD X60Y40VDD X65Y40VDD 25mOhm
L_X60Y40VDD_X70Y40VDD X65Y40VDD X70Y40VDD 2.91e-06nH
R_X60Y40VSS_X70Y40VSS X60Y40VSS X65Y40VSS 25mOhm
L_X60Y40VSS_X70Y40VSS X65Y40VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X80Y40VDD X70Y40VDD X75Y40VDD 25mOhm
L_X70Y40VDD_X80Y40VDD X75Y40VDD X80Y40VDD 2.91e-06nH
R_X70Y40VSS_X80Y40VSS X70Y40VSS X75Y40VSS 25mOhm
L_X70Y40VSS_X80Y40VSS X75Y40VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X90Y40VDD X80Y40VDD X85Y40VDD 25mOhm
L_X80Y40VDD_X90Y40VDD X85Y40VDD X90Y40VDD 2.91e-06nH
R_X80Y40VSS_X90Y40VSS X80Y40VSS X85Y40VSS 25mOhm
L_X80Y40VSS_X90Y40VSS X85Y40VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X100Y40VDD X90Y40VDD X95Y40VDD 25mOhm
L_X90Y40VDD_X100Y40VDD X95Y40VDD X100Y40VDD 2.91e-06nH
R_X90Y40VSS_X100Y40VSS X90Y40VSS X95Y40VSS 25mOhm
L_X90Y40VSS_X100Y40VSS X95Y40VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X110Y40VDD X100Y40VDD X105Y40VDD 25mOhm
L_X100Y40VDD_X110Y40VDD X105Y40VDD X110Y40VDD 2.91e-06nH
R_X100Y40VSS_X110Y40VSS X100Y40VSS X105Y40VSS 25mOhm
L_X100Y40VSS_X110Y40VSS X105Y40VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X120Y40VDD X110Y40VDD X115Y40VDD 25mOhm
L_X110Y40VDD_X120Y40VDD X115Y40VDD X120Y40VDD 2.91e-06nH
R_X110Y40VSS_X120Y40VSS X110Y40VSS X115Y40VSS 25mOhm
L_X110Y40VSS_X120Y40VSS X115Y40VSS X120Y40VSS 2.91e-06nH
R_X10Y50VDD_X20Y50VDD X10Y50VDD X15Y50VDD 25mOhm
L_X10Y50VDD_X20Y50VDD X15Y50VDD X20Y50VDD 2.91e-06nH
R_X10Y50VSS_X20Y50VSS X10Y50VSS X15Y50VSS 25mOhm
L_X10Y50VSS_X20Y50VSS X15Y50VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X30Y50VDD X20Y50VDD X25Y50VDD 25mOhm
L_X20Y50VDD_X30Y50VDD X25Y50VDD X30Y50VDD 2.91e-06nH
R_X20Y50VSS_X30Y50VSS X20Y50VSS X25Y50VSS 25mOhm
L_X20Y50VSS_X30Y50VSS X25Y50VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X40Y50VDD X30Y50VDD X35Y50VDD 25mOhm
L_X30Y50VDD_X40Y50VDD X35Y50VDD X40Y50VDD 2.91e-06nH
R_X30Y50VSS_X40Y50VSS X30Y50VSS X35Y50VSS 25mOhm
L_X30Y50VSS_X40Y50VSS X35Y50VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X50Y50VDD X40Y50VDD X45Y50VDD 25mOhm
L_X40Y50VDD_X50Y50VDD X45Y50VDD X50Y50VDD 2.91e-06nH
R_X40Y50VSS_X50Y50VSS X40Y50VSS X45Y50VSS 25mOhm
L_X40Y50VSS_X50Y50VSS X45Y50VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X60Y50VDD X50Y50VDD X55Y50VDD 25mOhm
L_X50Y50VDD_X60Y50VDD X55Y50VDD X60Y50VDD 2.91e-06nH
R_X50Y50VSS_X60Y50VSS X50Y50VSS X55Y50VSS 25mOhm
L_X50Y50VSS_X60Y50VSS X55Y50VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X70Y50VDD X60Y50VDD X65Y50VDD 25mOhm
L_X60Y50VDD_X70Y50VDD X65Y50VDD X70Y50VDD 2.91e-06nH
R_X60Y50VSS_X70Y50VSS X60Y50VSS X65Y50VSS 25mOhm
L_X60Y50VSS_X70Y50VSS X65Y50VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X80Y50VDD X70Y50VDD X75Y50VDD 25mOhm
L_X70Y50VDD_X80Y50VDD X75Y50VDD X80Y50VDD 2.91e-06nH
R_X70Y50VSS_X80Y50VSS X70Y50VSS X75Y50VSS 25mOhm
L_X70Y50VSS_X80Y50VSS X75Y50VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X90Y50VDD X80Y50VDD X85Y50VDD 25mOhm
L_X80Y50VDD_X90Y50VDD X85Y50VDD X90Y50VDD 2.91e-06nH
R_X80Y50VSS_X90Y50VSS X80Y50VSS X85Y50VSS 25mOhm
L_X80Y50VSS_X90Y50VSS X85Y50VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X100Y50VDD X90Y50VDD X95Y50VDD 25mOhm
L_X90Y50VDD_X100Y50VDD X95Y50VDD X100Y50VDD 2.91e-06nH
R_X90Y50VSS_X100Y50VSS X90Y50VSS X95Y50VSS 25mOhm
L_X90Y50VSS_X100Y50VSS X95Y50VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X110Y50VDD X100Y50VDD X105Y50VDD 25mOhm
L_X100Y50VDD_X110Y50VDD X105Y50VDD X110Y50VDD 2.91e-06nH
R_X100Y50VSS_X110Y50VSS X100Y50VSS X105Y50VSS 25mOhm
L_X100Y50VSS_X110Y50VSS X105Y50VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X120Y50VDD X110Y50VDD X115Y50VDD 25mOhm
L_X110Y50VDD_X120Y50VDD X115Y50VDD X120Y50VDD 2.91e-06nH
R_X110Y50VSS_X120Y50VSS X110Y50VSS X115Y50VSS 25mOhm
L_X110Y50VSS_X120Y50VSS X115Y50VSS X120Y50VSS 2.91e-06nH
R_X10Y60VDD_X20Y60VDD X10Y60VDD X15Y60VDD 25mOhm
L_X10Y60VDD_X20Y60VDD X15Y60VDD X20Y60VDD 2.91e-06nH
R_X10Y60VSS_X20Y60VSS X10Y60VSS X15Y60VSS 25mOhm
L_X10Y60VSS_X20Y60VSS X15Y60VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X30Y60VDD X20Y60VDD X25Y60VDD 25mOhm
L_X20Y60VDD_X30Y60VDD X25Y60VDD X30Y60VDD 2.91e-06nH
R_X20Y60VSS_X30Y60VSS X20Y60VSS X25Y60VSS 25mOhm
L_X20Y60VSS_X30Y60VSS X25Y60VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X40Y60VDD X30Y60VDD X35Y60VDD 25mOhm
L_X30Y60VDD_X40Y60VDD X35Y60VDD X40Y60VDD 2.91e-06nH
R_X30Y60VSS_X40Y60VSS X30Y60VSS X35Y60VSS 25mOhm
L_X30Y60VSS_X40Y60VSS X35Y60VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X50Y60VDD X40Y60VDD X45Y60VDD 25mOhm
L_X40Y60VDD_X50Y60VDD X45Y60VDD X50Y60VDD 2.91e-06nH
R_X40Y60VSS_X50Y60VSS X40Y60VSS X45Y60VSS 25mOhm
L_X40Y60VSS_X50Y60VSS X45Y60VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X60Y60VDD X50Y60VDD X55Y60VDD 25mOhm
L_X50Y60VDD_X60Y60VDD X55Y60VDD X60Y60VDD 2.91e-06nH
R_X50Y60VSS_X60Y60VSS X50Y60VSS X55Y60VSS 25mOhm
L_X50Y60VSS_X60Y60VSS X55Y60VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X70Y60VDD X60Y60VDD X65Y60VDD 25mOhm
L_X60Y60VDD_X70Y60VDD X65Y60VDD X70Y60VDD 2.91e-06nH
R_X60Y60VSS_X70Y60VSS X60Y60VSS X65Y60VSS 25mOhm
L_X60Y60VSS_X70Y60VSS X65Y60VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X80Y60VDD X70Y60VDD X75Y60VDD 25mOhm
L_X70Y60VDD_X80Y60VDD X75Y60VDD X80Y60VDD 2.91e-06nH
R_X70Y60VSS_X80Y60VSS X70Y60VSS X75Y60VSS 25mOhm
L_X70Y60VSS_X80Y60VSS X75Y60VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X90Y60VDD X80Y60VDD X85Y60VDD 25mOhm
L_X80Y60VDD_X90Y60VDD X85Y60VDD X90Y60VDD 2.91e-06nH
R_X80Y60VSS_X90Y60VSS X80Y60VSS X85Y60VSS 25mOhm
L_X80Y60VSS_X90Y60VSS X85Y60VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X100Y60VDD X90Y60VDD X95Y60VDD 25mOhm
L_X90Y60VDD_X100Y60VDD X95Y60VDD X100Y60VDD 2.91e-06nH
R_X90Y60VSS_X100Y60VSS X90Y60VSS X95Y60VSS 25mOhm
L_X90Y60VSS_X100Y60VSS X95Y60VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X110Y60VDD X100Y60VDD X105Y60VDD 25mOhm
L_X100Y60VDD_X110Y60VDD X105Y60VDD X110Y60VDD 2.91e-06nH
R_X100Y60VSS_X110Y60VSS X100Y60VSS X105Y60VSS 25mOhm
L_X100Y60VSS_X110Y60VSS X105Y60VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X120Y60VDD X110Y60VDD X115Y60VDD 25mOhm
L_X110Y60VDD_X120Y60VDD X115Y60VDD X120Y60VDD 2.91e-06nH
R_X110Y60VSS_X120Y60VSS X110Y60VSS X115Y60VSS 25mOhm
L_X110Y60VSS_X120Y60VSS X115Y60VSS X120Y60VSS 2.91e-06nH
R_X10Y70VDD_X20Y70VDD X10Y70VDD X15Y70VDD 25mOhm
L_X10Y70VDD_X20Y70VDD X15Y70VDD X20Y70VDD 2.91e-06nH
R_X10Y70VSS_X20Y70VSS X10Y70VSS X15Y70VSS 25mOhm
L_X10Y70VSS_X20Y70VSS X15Y70VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X30Y70VDD X20Y70VDD X25Y70VDD 25mOhm
L_X20Y70VDD_X30Y70VDD X25Y70VDD X30Y70VDD 2.91e-06nH
R_X20Y70VSS_X30Y70VSS X20Y70VSS X25Y70VSS 25mOhm
L_X20Y70VSS_X30Y70VSS X25Y70VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X40Y70VDD X30Y70VDD X35Y70VDD 25mOhm
L_X30Y70VDD_X40Y70VDD X35Y70VDD X40Y70VDD 2.91e-06nH
R_X30Y70VSS_X40Y70VSS X30Y70VSS X35Y70VSS 25mOhm
L_X30Y70VSS_X40Y70VSS X35Y70VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X50Y70VDD X40Y70VDD X45Y70VDD 25mOhm
L_X40Y70VDD_X50Y70VDD X45Y70VDD X50Y70VDD 2.91e-06nH
R_X40Y70VSS_X50Y70VSS X40Y70VSS X45Y70VSS 25mOhm
L_X40Y70VSS_X50Y70VSS X45Y70VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X60Y70VDD X50Y70VDD X55Y70VDD 25mOhm
L_X50Y70VDD_X60Y70VDD X55Y70VDD X60Y70VDD 2.91e-06nH
R_X50Y70VSS_X60Y70VSS X50Y70VSS X55Y70VSS 25mOhm
L_X50Y70VSS_X60Y70VSS X55Y70VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X70Y70VDD X60Y70VDD X65Y70VDD 25mOhm
L_X60Y70VDD_X70Y70VDD X65Y70VDD X70Y70VDD 2.91e-06nH
R_X60Y70VSS_X70Y70VSS X60Y70VSS X65Y70VSS 25mOhm
L_X60Y70VSS_X70Y70VSS X65Y70VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X80Y70VDD X70Y70VDD X75Y70VDD 25mOhm
L_X70Y70VDD_X80Y70VDD X75Y70VDD X80Y70VDD 2.91e-06nH
R_X70Y70VSS_X80Y70VSS X70Y70VSS X75Y70VSS 25mOhm
L_X70Y70VSS_X80Y70VSS X75Y70VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X90Y70VDD X80Y70VDD X85Y70VDD 25mOhm
L_X80Y70VDD_X90Y70VDD X85Y70VDD X90Y70VDD 2.91e-06nH
R_X80Y70VSS_X90Y70VSS X80Y70VSS X85Y70VSS 25mOhm
L_X80Y70VSS_X90Y70VSS X85Y70VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X100Y70VDD X90Y70VDD X95Y70VDD 25mOhm
L_X90Y70VDD_X100Y70VDD X95Y70VDD X100Y70VDD 2.91e-06nH
R_X90Y70VSS_X100Y70VSS X90Y70VSS X95Y70VSS 25mOhm
L_X90Y70VSS_X100Y70VSS X95Y70VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X110Y70VDD X100Y70VDD X105Y70VDD 25mOhm
L_X100Y70VDD_X110Y70VDD X105Y70VDD X110Y70VDD 2.91e-06nH
R_X100Y70VSS_X110Y70VSS X100Y70VSS X105Y70VSS 25mOhm
L_X100Y70VSS_X110Y70VSS X105Y70VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X120Y70VDD X110Y70VDD X115Y70VDD 25mOhm
L_X110Y70VDD_X120Y70VDD X115Y70VDD X120Y70VDD 2.91e-06nH
R_X110Y70VSS_X120Y70VSS X110Y70VSS X115Y70VSS 25mOhm
L_X110Y70VSS_X120Y70VSS X115Y70VSS X120Y70VSS 2.91e-06nH
R_X10Y80VDD_X20Y80VDD X10Y80VDD X15Y80VDD 25mOhm
L_X10Y80VDD_X20Y80VDD X15Y80VDD X20Y80VDD 2.91e-06nH
R_X10Y80VSS_X20Y80VSS X10Y80VSS X15Y80VSS 25mOhm
L_X10Y80VSS_X20Y80VSS X15Y80VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X30Y80VDD X20Y80VDD X25Y80VDD 25mOhm
L_X20Y80VDD_X30Y80VDD X25Y80VDD X30Y80VDD 2.91e-06nH
R_X20Y80VSS_X30Y80VSS X20Y80VSS X25Y80VSS 25mOhm
L_X20Y80VSS_X30Y80VSS X25Y80VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X40Y80VDD X30Y80VDD X35Y80VDD 25mOhm
L_X30Y80VDD_X40Y80VDD X35Y80VDD X40Y80VDD 2.91e-06nH
R_X30Y80VSS_X40Y80VSS X30Y80VSS X35Y80VSS 25mOhm
L_X30Y80VSS_X40Y80VSS X35Y80VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X50Y80VDD X40Y80VDD X45Y80VDD 25mOhm
L_X40Y80VDD_X50Y80VDD X45Y80VDD X50Y80VDD 2.91e-06nH
R_X40Y80VSS_X50Y80VSS X40Y80VSS X45Y80VSS 25mOhm
L_X40Y80VSS_X50Y80VSS X45Y80VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X60Y80VDD X50Y80VDD X55Y80VDD 25mOhm
L_X50Y80VDD_X60Y80VDD X55Y80VDD X60Y80VDD 2.91e-06nH
R_X50Y80VSS_X60Y80VSS X50Y80VSS X55Y80VSS 25mOhm
L_X50Y80VSS_X60Y80VSS X55Y80VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X70Y80VDD X60Y80VDD X65Y80VDD 25mOhm
L_X60Y80VDD_X70Y80VDD X65Y80VDD X70Y80VDD 2.91e-06nH
R_X60Y80VSS_X70Y80VSS X60Y80VSS X65Y80VSS 25mOhm
L_X60Y80VSS_X70Y80VSS X65Y80VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X80Y80VDD X70Y80VDD X75Y80VDD 25mOhm
L_X70Y80VDD_X80Y80VDD X75Y80VDD X80Y80VDD 2.91e-06nH
R_X70Y80VSS_X80Y80VSS X70Y80VSS X75Y80VSS 25mOhm
L_X70Y80VSS_X80Y80VSS X75Y80VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X90Y80VDD X80Y80VDD X85Y80VDD 25mOhm
L_X80Y80VDD_X90Y80VDD X85Y80VDD X90Y80VDD 2.91e-06nH
R_X80Y80VSS_X90Y80VSS X80Y80VSS X85Y80VSS 25mOhm
L_X80Y80VSS_X90Y80VSS X85Y80VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X100Y80VDD X90Y80VDD X95Y80VDD 25mOhm
L_X90Y80VDD_X100Y80VDD X95Y80VDD X100Y80VDD 2.91e-06nH
R_X90Y80VSS_X100Y80VSS X90Y80VSS X95Y80VSS 25mOhm
L_X90Y80VSS_X100Y80VSS X95Y80VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X110Y80VDD X100Y80VDD X105Y80VDD 25mOhm
L_X100Y80VDD_X110Y80VDD X105Y80VDD X110Y80VDD 2.91e-06nH
R_X100Y80VSS_X110Y80VSS X100Y80VSS X105Y80VSS 25mOhm
L_X100Y80VSS_X110Y80VSS X105Y80VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X120Y80VDD X110Y80VDD X115Y80VDD 25mOhm
L_X110Y80VDD_X120Y80VDD X115Y80VDD X120Y80VDD 2.91e-06nH
R_X110Y80VSS_X120Y80VSS X110Y80VSS X115Y80VSS 25mOhm
L_X110Y80VSS_X120Y80VSS X115Y80VSS X120Y80VSS 2.91e-06nH
R_X10Y90VDD_X20Y90VDD X10Y90VDD X15Y90VDD 25mOhm
L_X10Y90VDD_X20Y90VDD X15Y90VDD X20Y90VDD 2.91e-06nH
R_X10Y90VSS_X20Y90VSS X10Y90VSS X15Y90VSS 25mOhm
L_X10Y90VSS_X20Y90VSS X15Y90VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X30Y90VDD X20Y90VDD X25Y90VDD 25mOhm
L_X20Y90VDD_X30Y90VDD X25Y90VDD X30Y90VDD 2.91e-06nH
R_X20Y90VSS_X30Y90VSS X20Y90VSS X25Y90VSS 25mOhm
L_X20Y90VSS_X30Y90VSS X25Y90VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X40Y90VDD X30Y90VDD X35Y90VDD 25mOhm
L_X30Y90VDD_X40Y90VDD X35Y90VDD X40Y90VDD 2.91e-06nH
R_X30Y90VSS_X40Y90VSS X30Y90VSS X35Y90VSS 25mOhm
L_X30Y90VSS_X40Y90VSS X35Y90VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X50Y90VDD X40Y90VDD X45Y90VDD 25mOhm
L_X40Y90VDD_X50Y90VDD X45Y90VDD X50Y90VDD 2.91e-06nH
R_X40Y90VSS_X50Y90VSS X40Y90VSS X45Y90VSS 25mOhm
L_X40Y90VSS_X50Y90VSS X45Y90VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X60Y90VDD X50Y90VDD X55Y90VDD 25mOhm
L_X50Y90VDD_X60Y90VDD X55Y90VDD X60Y90VDD 2.91e-06nH
R_X50Y90VSS_X60Y90VSS X50Y90VSS X55Y90VSS 25mOhm
L_X50Y90VSS_X60Y90VSS X55Y90VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X70Y90VDD X60Y90VDD X65Y90VDD 25mOhm
L_X60Y90VDD_X70Y90VDD X65Y90VDD X70Y90VDD 2.91e-06nH
R_X60Y90VSS_X70Y90VSS X60Y90VSS X65Y90VSS 25mOhm
L_X60Y90VSS_X70Y90VSS X65Y90VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X80Y90VDD X70Y90VDD X75Y90VDD 25mOhm
L_X70Y90VDD_X80Y90VDD X75Y90VDD X80Y90VDD 2.91e-06nH
R_X70Y90VSS_X80Y90VSS X70Y90VSS X75Y90VSS 25mOhm
L_X70Y90VSS_X80Y90VSS X75Y90VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X90Y90VDD X80Y90VDD X85Y90VDD 25mOhm
L_X80Y90VDD_X90Y90VDD X85Y90VDD X90Y90VDD 2.91e-06nH
R_X80Y90VSS_X90Y90VSS X80Y90VSS X85Y90VSS 25mOhm
L_X80Y90VSS_X90Y90VSS X85Y90VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X100Y90VDD X90Y90VDD X95Y90VDD 25mOhm
L_X90Y90VDD_X100Y90VDD X95Y90VDD X100Y90VDD 2.91e-06nH
R_X90Y90VSS_X100Y90VSS X90Y90VSS X95Y90VSS 25mOhm
L_X90Y90VSS_X100Y90VSS X95Y90VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X110Y90VDD X100Y90VDD X105Y90VDD 25mOhm
L_X100Y90VDD_X110Y90VDD X105Y90VDD X110Y90VDD 2.91e-06nH
R_X100Y90VSS_X110Y90VSS X100Y90VSS X105Y90VSS 25mOhm
L_X100Y90VSS_X110Y90VSS X105Y90VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X120Y90VDD X110Y90VDD X115Y90VDD 25mOhm
L_X110Y90VDD_X120Y90VDD X115Y90VDD X120Y90VDD 2.91e-06nH
R_X110Y90VSS_X120Y90VSS X110Y90VSS X115Y90VSS 25mOhm
L_X110Y90VSS_X120Y90VSS X115Y90VSS X120Y90VSS 2.91e-06nH
R_X10Y100VDD_X20Y100VDD X10Y100VDD X15Y100VDD 25mOhm
L_X10Y100VDD_X20Y100VDD X15Y100VDD X20Y100VDD 2.91e-06nH
R_X10Y100VSS_X20Y100VSS X10Y100VSS X15Y100VSS 25mOhm
L_X10Y100VSS_X20Y100VSS X15Y100VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X30Y100VDD X20Y100VDD X25Y100VDD 25mOhm
L_X20Y100VDD_X30Y100VDD X25Y100VDD X30Y100VDD 2.91e-06nH
R_X20Y100VSS_X30Y100VSS X20Y100VSS X25Y100VSS 25mOhm
L_X20Y100VSS_X30Y100VSS X25Y100VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X40Y100VDD X30Y100VDD X35Y100VDD 25mOhm
L_X30Y100VDD_X40Y100VDD X35Y100VDD X40Y100VDD 2.91e-06nH
R_X30Y100VSS_X40Y100VSS X30Y100VSS X35Y100VSS 25mOhm
L_X30Y100VSS_X40Y100VSS X35Y100VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X50Y100VDD X40Y100VDD X45Y100VDD 25mOhm
L_X40Y100VDD_X50Y100VDD X45Y100VDD X50Y100VDD 2.91e-06nH
R_X40Y100VSS_X50Y100VSS X40Y100VSS X45Y100VSS 25mOhm
L_X40Y100VSS_X50Y100VSS X45Y100VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X60Y100VDD X50Y100VDD X55Y100VDD 25mOhm
L_X50Y100VDD_X60Y100VDD X55Y100VDD X60Y100VDD 2.91e-06nH
R_X50Y100VSS_X60Y100VSS X50Y100VSS X55Y100VSS 25mOhm
L_X50Y100VSS_X60Y100VSS X55Y100VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X70Y100VDD X60Y100VDD X65Y100VDD 25mOhm
L_X60Y100VDD_X70Y100VDD X65Y100VDD X70Y100VDD 2.91e-06nH
R_X60Y100VSS_X70Y100VSS X60Y100VSS X65Y100VSS 25mOhm
L_X60Y100VSS_X70Y100VSS X65Y100VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X80Y100VDD X70Y100VDD X75Y100VDD 25mOhm
L_X70Y100VDD_X80Y100VDD X75Y100VDD X80Y100VDD 2.91e-06nH
R_X70Y100VSS_X80Y100VSS X70Y100VSS X75Y100VSS 25mOhm
L_X70Y100VSS_X80Y100VSS X75Y100VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X90Y100VDD X80Y100VDD X85Y100VDD 25mOhm
L_X80Y100VDD_X90Y100VDD X85Y100VDD X90Y100VDD 2.91e-06nH
R_X80Y100VSS_X90Y100VSS X80Y100VSS X85Y100VSS 25mOhm
L_X80Y100VSS_X90Y100VSS X85Y100VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X100Y100VDD X90Y100VDD X95Y100VDD 25mOhm
L_X90Y100VDD_X100Y100VDD X95Y100VDD X100Y100VDD 2.91e-06nH
R_X90Y100VSS_X100Y100VSS X90Y100VSS X95Y100VSS 25mOhm
L_X90Y100VSS_X100Y100VSS X95Y100VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X110Y100VDD X100Y100VDD X105Y100VDD 25mOhm
L_X100Y100VDD_X110Y100VDD X105Y100VDD X110Y100VDD 2.91e-06nH
R_X100Y100VSS_X110Y100VSS X100Y100VSS X105Y100VSS 25mOhm
L_X100Y100VSS_X110Y100VSS X105Y100VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X120Y100VDD X110Y100VDD X115Y100VDD 25mOhm
L_X110Y100VDD_X120Y100VDD X115Y100VDD X120Y100VDD 2.91e-06nH
R_X110Y100VSS_X120Y100VSS X110Y100VSS X115Y100VSS 25mOhm
L_X110Y100VSS_X120Y100VSS X115Y100VSS X120Y100VSS 2.91e-06nH
R_X10Y110VDD_X20Y110VDD X10Y110VDD X15Y110VDD 25mOhm
L_X10Y110VDD_X20Y110VDD X15Y110VDD X20Y110VDD 2.91e-06nH
R_X10Y110VSS_X20Y110VSS X10Y110VSS X15Y110VSS 25mOhm
L_X10Y110VSS_X20Y110VSS X15Y110VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X30Y110VDD X20Y110VDD X25Y110VDD 25mOhm
L_X20Y110VDD_X30Y110VDD X25Y110VDD X30Y110VDD 2.91e-06nH
R_X20Y110VSS_X30Y110VSS X20Y110VSS X25Y110VSS 25mOhm
L_X20Y110VSS_X30Y110VSS X25Y110VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X40Y110VDD X30Y110VDD X35Y110VDD 25mOhm
L_X30Y110VDD_X40Y110VDD X35Y110VDD X40Y110VDD 2.91e-06nH
R_X30Y110VSS_X40Y110VSS X30Y110VSS X35Y110VSS 25mOhm
L_X30Y110VSS_X40Y110VSS X35Y110VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X50Y110VDD X40Y110VDD X45Y110VDD 25mOhm
L_X40Y110VDD_X50Y110VDD X45Y110VDD X50Y110VDD 2.91e-06nH
R_X40Y110VSS_X50Y110VSS X40Y110VSS X45Y110VSS 25mOhm
L_X40Y110VSS_X50Y110VSS X45Y110VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X60Y110VDD X50Y110VDD X55Y110VDD 25mOhm
L_X50Y110VDD_X60Y110VDD X55Y110VDD X60Y110VDD 2.91e-06nH
R_X50Y110VSS_X60Y110VSS X50Y110VSS X55Y110VSS 25mOhm
L_X50Y110VSS_X60Y110VSS X55Y110VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X70Y110VDD X60Y110VDD X65Y110VDD 25mOhm
L_X60Y110VDD_X70Y110VDD X65Y110VDD X70Y110VDD 2.91e-06nH
R_X60Y110VSS_X70Y110VSS X60Y110VSS X65Y110VSS 25mOhm
L_X60Y110VSS_X70Y110VSS X65Y110VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X80Y110VDD X70Y110VDD X75Y110VDD 25mOhm
L_X70Y110VDD_X80Y110VDD X75Y110VDD X80Y110VDD 2.91e-06nH
R_X70Y110VSS_X80Y110VSS X70Y110VSS X75Y110VSS 25mOhm
L_X70Y110VSS_X80Y110VSS X75Y110VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X90Y110VDD X80Y110VDD X85Y110VDD 25mOhm
L_X80Y110VDD_X90Y110VDD X85Y110VDD X90Y110VDD 2.91e-06nH
R_X80Y110VSS_X90Y110VSS X80Y110VSS X85Y110VSS 25mOhm
L_X80Y110VSS_X90Y110VSS X85Y110VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X100Y110VDD X90Y110VDD X95Y110VDD 25mOhm
L_X90Y110VDD_X100Y110VDD X95Y110VDD X100Y110VDD 2.91e-06nH
R_X90Y110VSS_X100Y110VSS X90Y110VSS X95Y110VSS 25mOhm
L_X90Y110VSS_X100Y110VSS X95Y110VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X110Y110VDD X100Y110VDD X105Y110VDD 25mOhm
L_X100Y110VDD_X110Y110VDD X105Y110VDD X110Y110VDD 2.91e-06nH
R_X100Y110VSS_X110Y110VSS X100Y110VSS X105Y110VSS 25mOhm
L_X100Y110VSS_X110Y110VSS X105Y110VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X120Y110VDD X110Y110VDD X115Y110VDD 25mOhm
L_X110Y110VDD_X120Y110VDD X115Y110VDD X120Y110VDD 2.91e-06nH
R_X110Y110VSS_X120Y110VSS X110Y110VSS X115Y110VSS 25mOhm
L_X110Y110VSS_X120Y110VSS X115Y110VSS X120Y110VSS 2.91e-06nH
R_X10Y120VDD_X20Y120VDD X10Y120VDD X15Y120VDD 25mOhm
L_X10Y120VDD_X20Y120VDD X15Y120VDD X20Y120VDD 2.91e-06nH
R_X10Y120VSS_X20Y120VSS X10Y120VSS X15Y120VSS 25mOhm
L_X10Y120VSS_X20Y120VSS X15Y120VSS X20Y120VSS 2.91e-06nH
R_X20Y120VDD_X30Y120VDD X20Y120VDD X25Y120VDD 25mOhm
L_X20Y120VDD_X30Y120VDD X25Y120VDD X30Y120VDD 2.91e-06nH
R_X20Y120VSS_X30Y120VSS X20Y120VSS X25Y120VSS 25mOhm
L_X20Y120VSS_X30Y120VSS X25Y120VSS X30Y120VSS 2.91e-06nH
R_X30Y120VDD_X40Y120VDD X30Y120VDD X35Y120VDD 25mOhm
L_X30Y120VDD_X40Y120VDD X35Y120VDD X40Y120VDD 2.91e-06nH
R_X30Y120VSS_X40Y120VSS X30Y120VSS X35Y120VSS 25mOhm
L_X30Y120VSS_X40Y120VSS X35Y120VSS X40Y120VSS 2.91e-06nH
R_X40Y120VDD_X50Y120VDD X40Y120VDD X45Y120VDD 25mOhm
L_X40Y120VDD_X50Y120VDD X45Y120VDD X50Y120VDD 2.91e-06nH
R_X40Y120VSS_X50Y120VSS X40Y120VSS X45Y120VSS 25mOhm
L_X40Y120VSS_X50Y120VSS X45Y120VSS X50Y120VSS 2.91e-06nH
R_X50Y120VDD_X60Y120VDD X50Y120VDD X55Y120VDD 25mOhm
L_X50Y120VDD_X60Y120VDD X55Y120VDD X60Y120VDD 2.91e-06nH
R_X50Y120VSS_X60Y120VSS X50Y120VSS X55Y120VSS 25mOhm
L_X50Y120VSS_X60Y120VSS X55Y120VSS X60Y120VSS 2.91e-06nH
R_X60Y120VDD_X70Y120VDD X60Y120VDD X65Y120VDD 25mOhm
L_X60Y120VDD_X70Y120VDD X65Y120VDD X70Y120VDD 2.91e-06nH
R_X60Y120VSS_X70Y120VSS X60Y120VSS X65Y120VSS 25mOhm
L_X60Y120VSS_X70Y120VSS X65Y120VSS X70Y120VSS 2.91e-06nH
R_X70Y120VDD_X80Y120VDD X70Y120VDD X75Y120VDD 25mOhm
L_X70Y120VDD_X80Y120VDD X75Y120VDD X80Y120VDD 2.91e-06nH
R_X70Y120VSS_X80Y120VSS X70Y120VSS X75Y120VSS 25mOhm
L_X70Y120VSS_X80Y120VSS X75Y120VSS X80Y120VSS 2.91e-06nH
R_X80Y120VDD_X90Y120VDD X80Y120VDD X85Y120VDD 25mOhm
L_X80Y120VDD_X90Y120VDD X85Y120VDD X90Y120VDD 2.91e-06nH
R_X80Y120VSS_X90Y120VSS X80Y120VSS X85Y120VSS 25mOhm
L_X80Y120VSS_X90Y120VSS X85Y120VSS X90Y120VSS 2.91e-06nH
R_X90Y120VDD_X100Y120VDD X90Y120VDD X95Y120VDD 25mOhm
L_X90Y120VDD_X100Y120VDD X95Y120VDD X100Y120VDD 2.91e-06nH
R_X90Y120VSS_X100Y120VSS X90Y120VSS X95Y120VSS 25mOhm
L_X90Y120VSS_X100Y120VSS X95Y120VSS X100Y120VSS 2.91e-06nH
R_X100Y120VDD_X110Y120VDD X100Y120VDD X105Y120VDD 25mOhm
L_X100Y120VDD_X110Y120VDD X105Y120VDD X110Y120VDD 2.91e-06nH
R_X100Y120VSS_X110Y120VSS X100Y120VSS X105Y120VSS 25mOhm
L_X100Y120VSS_X110Y120VSS X105Y120VSS X110Y120VSS 2.91e-06nH
R_X110Y120VDD_X120Y120VDD X110Y120VDD X115Y120VDD 25mOhm
L_X110Y120VDD_X120Y120VDD X115Y120VDD X120Y120VDD 2.91e-06nH
R_X110Y120VSS_X120Y120VSS X110Y120VSS X115Y120VSS 25mOhm
L_X110Y120VSS_X120Y120VSS X115Y120VSS X120Y120VSS 2.91e-06nH
R_X10Y10VDD_X10Y20VDD X10Y10VDD X10Y15VDD 25mOhm
L_X10Y10VDD_X10Y20VDD X10Y15VDD X10Y20VDD 2.91e-06nH
R_X10Y10VSS_X10Y20VSS X10Y10VSS X10Y15VSS 25mOhm
L_X10Y10VSS_X10Y20VSS X10Y15VSS X10Y20VSS 2.91e-06nH
R_X10Y20VDD_X10Y30VDD X10Y20VDD X10Y25VDD 25mOhm
L_X10Y20VDD_X10Y30VDD X10Y25VDD X10Y30VDD 2.91e-06nH
R_X10Y20VSS_X10Y30VSS X10Y20VSS X10Y25VSS 25mOhm
L_X10Y20VSS_X10Y30VSS X10Y25VSS X10Y30VSS 2.91e-06nH
R_X10Y30VDD_X10Y40VDD X10Y30VDD X10Y35VDD 25mOhm
L_X10Y30VDD_X10Y40VDD X10Y35VDD X10Y40VDD 2.91e-06nH
R_X10Y30VSS_X10Y40VSS X10Y30VSS X10Y35VSS 25mOhm
L_X10Y30VSS_X10Y40VSS X10Y35VSS X10Y40VSS 2.91e-06nH
R_X10Y40VDD_X10Y50VDD X10Y40VDD X10Y45VDD 25mOhm
L_X10Y40VDD_X10Y50VDD X10Y45VDD X10Y50VDD 2.91e-06nH
R_X10Y40VSS_X10Y50VSS X10Y40VSS X10Y45VSS 25mOhm
L_X10Y40VSS_X10Y50VSS X10Y45VSS X10Y50VSS 2.91e-06nH
R_X10Y50VDD_X10Y60VDD X10Y50VDD X10Y55VDD 25mOhm
L_X10Y50VDD_X10Y60VDD X10Y55VDD X10Y60VDD 2.91e-06nH
R_X10Y50VSS_X10Y60VSS X10Y50VSS X10Y55VSS 25mOhm
L_X10Y50VSS_X10Y60VSS X10Y55VSS X10Y60VSS 2.91e-06nH
R_X10Y60VDD_X10Y70VDD X10Y60VDD X10Y65VDD 25mOhm
L_X10Y60VDD_X10Y70VDD X10Y65VDD X10Y70VDD 2.91e-06nH
R_X10Y60VSS_X10Y70VSS X10Y60VSS X10Y65VSS 25mOhm
L_X10Y60VSS_X10Y70VSS X10Y65VSS X10Y70VSS 2.91e-06nH
R_X10Y70VDD_X10Y80VDD X10Y70VDD X10Y75VDD 25mOhm
L_X10Y70VDD_X10Y80VDD X10Y75VDD X10Y80VDD 2.91e-06nH
R_X10Y70VSS_X10Y80VSS X10Y70VSS X10Y75VSS 25mOhm
L_X10Y70VSS_X10Y80VSS X10Y75VSS X10Y80VSS 2.91e-06nH
R_X10Y80VDD_X10Y90VDD X10Y80VDD X10Y85VDD 25mOhm
L_X10Y80VDD_X10Y90VDD X10Y85VDD X10Y90VDD 2.91e-06nH
R_X10Y80VSS_X10Y90VSS X10Y80VSS X10Y85VSS 25mOhm
L_X10Y80VSS_X10Y90VSS X10Y85VSS X10Y90VSS 2.91e-06nH
R_X10Y90VDD_X10Y100VDD X10Y90VDD X10Y95VDD 25mOhm
L_X10Y90VDD_X10Y100VDD X10Y95VDD X10Y100VDD 2.91e-06nH
R_X10Y90VSS_X10Y100VSS X10Y90VSS X10Y95VSS 25mOhm
L_X10Y90VSS_X10Y100VSS X10Y95VSS X10Y100VSS 2.91e-06nH
R_X10Y100VDD_X10Y110VDD X10Y100VDD X10Y105VDD 25mOhm
L_X10Y100VDD_X10Y110VDD X10Y105VDD X10Y110VDD 2.91e-06nH
R_X10Y100VSS_X10Y110VSS X10Y100VSS X10Y105VSS 25mOhm
L_X10Y100VSS_X10Y110VSS X10Y105VSS X10Y110VSS 2.91e-06nH
R_X10Y110VDD_X10Y120VDD X10Y110VDD X10Y115VDD 25mOhm
L_X10Y110VDD_X10Y120VDD X10Y115VDD X10Y120VDD 2.91e-06nH
R_X10Y110VSS_X10Y120VSS X10Y110VSS X10Y115VSS 25mOhm
L_X10Y110VSS_X10Y120VSS X10Y115VSS X10Y120VSS 2.91e-06nH
R_X20Y10VDD_X20Y20VDD X20Y10VDD X20Y15VDD 25mOhm
L_X20Y10VDD_X20Y20VDD X20Y15VDD X20Y20VDD 2.91e-06nH
R_X20Y10VSS_X20Y20VSS X20Y10VSS X20Y15VSS 25mOhm
L_X20Y10VSS_X20Y20VSS X20Y15VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X20Y30VDD X20Y20VDD X20Y25VDD 25mOhm
L_X20Y20VDD_X20Y30VDD X20Y25VDD X20Y30VDD 2.91e-06nH
R_X20Y20VSS_X20Y30VSS X20Y20VSS X20Y25VSS 25mOhm
L_X20Y20VSS_X20Y30VSS X20Y25VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X20Y40VDD X20Y30VDD X20Y35VDD 25mOhm
L_X20Y30VDD_X20Y40VDD X20Y35VDD X20Y40VDD 2.91e-06nH
R_X20Y30VSS_X20Y40VSS X20Y30VSS X20Y35VSS 25mOhm
L_X20Y30VSS_X20Y40VSS X20Y35VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X20Y50VDD X20Y40VDD X20Y45VDD 25mOhm
L_X20Y40VDD_X20Y50VDD X20Y45VDD X20Y50VDD 2.91e-06nH
R_X20Y40VSS_X20Y50VSS X20Y40VSS X20Y45VSS 25mOhm
L_X20Y40VSS_X20Y50VSS X20Y45VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X20Y60VDD X20Y50VDD X20Y55VDD 25mOhm
L_X20Y50VDD_X20Y60VDD X20Y55VDD X20Y60VDD 2.91e-06nH
R_X20Y50VSS_X20Y60VSS X20Y50VSS X20Y55VSS 25mOhm
L_X20Y50VSS_X20Y60VSS X20Y55VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X20Y70VDD X20Y60VDD X20Y65VDD 25mOhm
L_X20Y60VDD_X20Y70VDD X20Y65VDD X20Y70VDD 2.91e-06nH
R_X20Y60VSS_X20Y70VSS X20Y60VSS X20Y65VSS 25mOhm
L_X20Y60VSS_X20Y70VSS X20Y65VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X20Y80VDD X20Y70VDD X20Y75VDD 25mOhm
L_X20Y70VDD_X20Y80VDD X20Y75VDD X20Y80VDD 2.91e-06nH
R_X20Y70VSS_X20Y80VSS X20Y70VSS X20Y75VSS 25mOhm
L_X20Y70VSS_X20Y80VSS X20Y75VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X20Y90VDD X20Y80VDD X20Y85VDD 25mOhm
L_X20Y80VDD_X20Y90VDD X20Y85VDD X20Y90VDD 2.91e-06nH
R_X20Y80VSS_X20Y90VSS X20Y80VSS X20Y85VSS 25mOhm
L_X20Y80VSS_X20Y90VSS X20Y85VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X20Y100VDD X20Y90VDD X20Y95VDD 25mOhm
L_X20Y90VDD_X20Y100VDD X20Y95VDD X20Y100VDD 2.91e-06nH
R_X20Y90VSS_X20Y100VSS X20Y90VSS X20Y95VSS 25mOhm
L_X20Y90VSS_X20Y100VSS X20Y95VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X20Y110VDD X20Y100VDD X20Y105VDD 25mOhm
L_X20Y100VDD_X20Y110VDD X20Y105VDD X20Y110VDD 2.91e-06nH
R_X20Y100VSS_X20Y110VSS X20Y100VSS X20Y105VSS 25mOhm
L_X20Y100VSS_X20Y110VSS X20Y105VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X20Y120VDD X20Y110VDD X20Y115VDD 25mOhm
L_X20Y110VDD_X20Y120VDD X20Y115VDD X20Y120VDD 2.91e-06nH
R_X20Y110VSS_X20Y120VSS X20Y110VSS X20Y115VSS 25mOhm
L_X20Y110VSS_X20Y120VSS X20Y115VSS X20Y120VSS 2.91e-06nH
R_X30Y10VDD_X30Y20VDD X30Y10VDD X30Y15VDD 25mOhm
L_X30Y10VDD_X30Y20VDD X30Y15VDD X30Y20VDD 2.91e-06nH
R_X30Y10VSS_X30Y20VSS X30Y10VSS X30Y15VSS 25mOhm
L_X30Y10VSS_X30Y20VSS X30Y15VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X30Y30VDD X30Y20VDD X30Y25VDD 25mOhm
L_X30Y20VDD_X30Y30VDD X30Y25VDD X30Y30VDD 2.91e-06nH
R_X30Y20VSS_X30Y30VSS X30Y20VSS X30Y25VSS 25mOhm
L_X30Y20VSS_X30Y30VSS X30Y25VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X30Y40VDD X30Y30VDD X30Y35VDD 25mOhm
L_X30Y30VDD_X30Y40VDD X30Y35VDD X30Y40VDD 2.91e-06nH
R_X30Y30VSS_X30Y40VSS X30Y30VSS X30Y35VSS 25mOhm
L_X30Y30VSS_X30Y40VSS X30Y35VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X30Y50VDD X30Y40VDD X30Y45VDD 25mOhm
L_X30Y40VDD_X30Y50VDD X30Y45VDD X30Y50VDD 2.91e-06nH
R_X30Y40VSS_X30Y50VSS X30Y40VSS X30Y45VSS 25mOhm
L_X30Y40VSS_X30Y50VSS X30Y45VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X30Y60VDD X30Y50VDD X30Y55VDD 25mOhm
L_X30Y50VDD_X30Y60VDD X30Y55VDD X30Y60VDD 2.91e-06nH
R_X30Y50VSS_X30Y60VSS X30Y50VSS X30Y55VSS 25mOhm
L_X30Y50VSS_X30Y60VSS X30Y55VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X30Y70VDD X30Y60VDD X30Y65VDD 25mOhm
L_X30Y60VDD_X30Y70VDD X30Y65VDD X30Y70VDD 2.91e-06nH
R_X30Y60VSS_X30Y70VSS X30Y60VSS X30Y65VSS 25mOhm
L_X30Y60VSS_X30Y70VSS X30Y65VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X30Y80VDD X30Y70VDD X30Y75VDD 25mOhm
L_X30Y70VDD_X30Y80VDD X30Y75VDD X30Y80VDD 2.91e-06nH
R_X30Y70VSS_X30Y80VSS X30Y70VSS X30Y75VSS 25mOhm
L_X30Y70VSS_X30Y80VSS X30Y75VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X30Y90VDD X30Y80VDD X30Y85VDD 25mOhm
L_X30Y80VDD_X30Y90VDD X30Y85VDD X30Y90VDD 2.91e-06nH
R_X30Y80VSS_X30Y90VSS X30Y80VSS X30Y85VSS 25mOhm
L_X30Y80VSS_X30Y90VSS X30Y85VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X30Y100VDD X30Y90VDD X30Y95VDD 25mOhm
L_X30Y90VDD_X30Y100VDD X30Y95VDD X30Y100VDD 2.91e-06nH
R_X30Y90VSS_X30Y100VSS X30Y90VSS X30Y95VSS 25mOhm
L_X30Y90VSS_X30Y100VSS X30Y95VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X30Y110VDD X30Y100VDD X30Y105VDD 25mOhm
L_X30Y100VDD_X30Y110VDD X30Y105VDD X30Y110VDD 2.91e-06nH
R_X30Y100VSS_X30Y110VSS X30Y100VSS X30Y105VSS 25mOhm
L_X30Y100VSS_X30Y110VSS X30Y105VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X30Y120VDD X30Y110VDD X30Y115VDD 25mOhm
L_X30Y110VDD_X30Y120VDD X30Y115VDD X30Y120VDD 2.91e-06nH
R_X30Y110VSS_X30Y120VSS X30Y110VSS X30Y115VSS 25mOhm
L_X30Y110VSS_X30Y120VSS X30Y115VSS X30Y120VSS 2.91e-06nH
R_X40Y10VDD_X40Y20VDD X40Y10VDD X40Y15VDD 25mOhm
L_X40Y10VDD_X40Y20VDD X40Y15VDD X40Y20VDD 2.91e-06nH
R_X40Y10VSS_X40Y20VSS X40Y10VSS X40Y15VSS 25mOhm
L_X40Y10VSS_X40Y20VSS X40Y15VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X40Y30VDD X40Y20VDD X40Y25VDD 25mOhm
L_X40Y20VDD_X40Y30VDD X40Y25VDD X40Y30VDD 2.91e-06nH
R_X40Y20VSS_X40Y30VSS X40Y20VSS X40Y25VSS 25mOhm
L_X40Y20VSS_X40Y30VSS X40Y25VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X40Y40VDD X40Y30VDD X40Y35VDD 25mOhm
L_X40Y30VDD_X40Y40VDD X40Y35VDD X40Y40VDD 2.91e-06nH
R_X40Y30VSS_X40Y40VSS X40Y30VSS X40Y35VSS 25mOhm
L_X40Y30VSS_X40Y40VSS X40Y35VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X40Y50VDD X40Y40VDD X40Y45VDD 25mOhm
L_X40Y40VDD_X40Y50VDD X40Y45VDD X40Y50VDD 2.91e-06nH
R_X40Y40VSS_X40Y50VSS X40Y40VSS X40Y45VSS 25mOhm
L_X40Y40VSS_X40Y50VSS X40Y45VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X40Y60VDD X40Y50VDD X40Y55VDD 25mOhm
L_X40Y50VDD_X40Y60VDD X40Y55VDD X40Y60VDD 2.91e-06nH
R_X40Y50VSS_X40Y60VSS X40Y50VSS X40Y55VSS 25mOhm
L_X40Y50VSS_X40Y60VSS X40Y55VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X40Y70VDD X40Y60VDD X40Y65VDD 25mOhm
L_X40Y60VDD_X40Y70VDD X40Y65VDD X40Y70VDD 2.91e-06nH
R_X40Y60VSS_X40Y70VSS X40Y60VSS X40Y65VSS 25mOhm
L_X40Y60VSS_X40Y70VSS X40Y65VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X40Y80VDD X40Y70VDD X40Y75VDD 25mOhm
L_X40Y70VDD_X40Y80VDD X40Y75VDD X40Y80VDD 2.91e-06nH
R_X40Y70VSS_X40Y80VSS X40Y70VSS X40Y75VSS 25mOhm
L_X40Y70VSS_X40Y80VSS X40Y75VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X40Y90VDD X40Y80VDD X40Y85VDD 25mOhm
L_X40Y80VDD_X40Y90VDD X40Y85VDD X40Y90VDD 2.91e-06nH
R_X40Y80VSS_X40Y90VSS X40Y80VSS X40Y85VSS 25mOhm
L_X40Y80VSS_X40Y90VSS X40Y85VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X40Y100VDD X40Y90VDD X40Y95VDD 25mOhm
L_X40Y90VDD_X40Y100VDD X40Y95VDD X40Y100VDD 2.91e-06nH
R_X40Y90VSS_X40Y100VSS X40Y90VSS X40Y95VSS 25mOhm
L_X40Y90VSS_X40Y100VSS X40Y95VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X40Y110VDD X40Y100VDD X40Y105VDD 25mOhm
L_X40Y100VDD_X40Y110VDD X40Y105VDD X40Y110VDD 2.91e-06nH
R_X40Y100VSS_X40Y110VSS X40Y100VSS X40Y105VSS 25mOhm
L_X40Y100VSS_X40Y110VSS X40Y105VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X40Y120VDD X40Y110VDD X40Y115VDD 25mOhm
L_X40Y110VDD_X40Y120VDD X40Y115VDD X40Y120VDD 2.91e-06nH
R_X40Y110VSS_X40Y120VSS X40Y110VSS X40Y115VSS 25mOhm
L_X40Y110VSS_X40Y120VSS X40Y115VSS X40Y120VSS 2.91e-06nH
R_X50Y10VDD_X50Y20VDD X50Y10VDD X50Y15VDD 25mOhm
L_X50Y10VDD_X50Y20VDD X50Y15VDD X50Y20VDD 2.91e-06nH
R_X50Y10VSS_X50Y20VSS X50Y10VSS X50Y15VSS 25mOhm
L_X50Y10VSS_X50Y20VSS X50Y15VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X50Y30VDD X50Y20VDD X50Y25VDD 25mOhm
L_X50Y20VDD_X50Y30VDD X50Y25VDD X50Y30VDD 2.91e-06nH
R_X50Y20VSS_X50Y30VSS X50Y20VSS X50Y25VSS 25mOhm
L_X50Y20VSS_X50Y30VSS X50Y25VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X50Y40VDD X50Y30VDD X50Y35VDD 25mOhm
L_X50Y30VDD_X50Y40VDD X50Y35VDD X50Y40VDD 2.91e-06nH
R_X50Y30VSS_X50Y40VSS X50Y30VSS X50Y35VSS 25mOhm
L_X50Y30VSS_X50Y40VSS X50Y35VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X50Y50VDD X50Y40VDD X50Y45VDD 25mOhm
L_X50Y40VDD_X50Y50VDD X50Y45VDD X50Y50VDD 2.91e-06nH
R_X50Y40VSS_X50Y50VSS X50Y40VSS X50Y45VSS 25mOhm
L_X50Y40VSS_X50Y50VSS X50Y45VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X50Y60VDD X50Y50VDD X50Y55VDD 25mOhm
L_X50Y50VDD_X50Y60VDD X50Y55VDD X50Y60VDD 2.91e-06nH
R_X50Y50VSS_X50Y60VSS X50Y50VSS X50Y55VSS 25mOhm
L_X50Y50VSS_X50Y60VSS X50Y55VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X50Y70VDD X50Y60VDD X50Y65VDD 25mOhm
L_X50Y60VDD_X50Y70VDD X50Y65VDD X50Y70VDD 2.91e-06nH
R_X50Y60VSS_X50Y70VSS X50Y60VSS X50Y65VSS 25mOhm
L_X50Y60VSS_X50Y70VSS X50Y65VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X50Y80VDD X50Y70VDD X50Y75VDD 25mOhm
L_X50Y70VDD_X50Y80VDD X50Y75VDD X50Y80VDD 2.91e-06nH
R_X50Y70VSS_X50Y80VSS X50Y70VSS X50Y75VSS 25mOhm
L_X50Y70VSS_X50Y80VSS X50Y75VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X50Y90VDD X50Y80VDD X50Y85VDD 25mOhm
L_X50Y80VDD_X50Y90VDD X50Y85VDD X50Y90VDD 2.91e-06nH
R_X50Y80VSS_X50Y90VSS X50Y80VSS X50Y85VSS 25mOhm
L_X50Y80VSS_X50Y90VSS X50Y85VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X50Y100VDD X50Y90VDD X50Y95VDD 25mOhm
L_X50Y90VDD_X50Y100VDD X50Y95VDD X50Y100VDD 2.91e-06nH
R_X50Y90VSS_X50Y100VSS X50Y90VSS X50Y95VSS 25mOhm
L_X50Y90VSS_X50Y100VSS X50Y95VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X50Y110VDD X50Y100VDD X50Y105VDD 25mOhm
L_X50Y100VDD_X50Y110VDD X50Y105VDD X50Y110VDD 2.91e-06nH
R_X50Y100VSS_X50Y110VSS X50Y100VSS X50Y105VSS 25mOhm
L_X50Y100VSS_X50Y110VSS X50Y105VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X50Y120VDD X50Y110VDD X50Y115VDD 25mOhm
L_X50Y110VDD_X50Y120VDD X50Y115VDD X50Y120VDD 2.91e-06nH
R_X50Y110VSS_X50Y120VSS X50Y110VSS X50Y115VSS 25mOhm
L_X50Y110VSS_X50Y120VSS X50Y115VSS X50Y120VSS 2.91e-06nH
R_X60Y10VDD_X60Y20VDD X60Y10VDD X60Y15VDD 25mOhm
L_X60Y10VDD_X60Y20VDD X60Y15VDD X60Y20VDD 2.91e-06nH
R_X60Y10VSS_X60Y20VSS X60Y10VSS X60Y15VSS 25mOhm
L_X60Y10VSS_X60Y20VSS X60Y15VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X60Y30VDD X60Y20VDD X60Y25VDD 25mOhm
L_X60Y20VDD_X60Y30VDD X60Y25VDD X60Y30VDD 2.91e-06nH
R_X60Y20VSS_X60Y30VSS X60Y20VSS X60Y25VSS 25mOhm
L_X60Y20VSS_X60Y30VSS X60Y25VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X60Y40VDD X60Y30VDD X60Y35VDD 25mOhm
L_X60Y30VDD_X60Y40VDD X60Y35VDD X60Y40VDD 2.91e-06nH
R_X60Y30VSS_X60Y40VSS X60Y30VSS X60Y35VSS 25mOhm
L_X60Y30VSS_X60Y40VSS X60Y35VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X60Y50VDD X60Y40VDD X60Y45VDD 25mOhm
L_X60Y40VDD_X60Y50VDD X60Y45VDD X60Y50VDD 2.91e-06nH
R_X60Y40VSS_X60Y50VSS X60Y40VSS X60Y45VSS 25mOhm
L_X60Y40VSS_X60Y50VSS X60Y45VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X60Y60VDD X60Y50VDD X60Y55VDD 25mOhm
L_X60Y50VDD_X60Y60VDD X60Y55VDD X60Y60VDD 2.91e-06nH
R_X60Y50VSS_X60Y60VSS X60Y50VSS X60Y55VSS 25mOhm
L_X60Y50VSS_X60Y60VSS X60Y55VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X60Y70VDD X60Y60VDD X60Y65VDD 25mOhm
L_X60Y60VDD_X60Y70VDD X60Y65VDD X60Y70VDD 2.91e-06nH
R_X60Y60VSS_X60Y70VSS X60Y60VSS X60Y65VSS 25mOhm
L_X60Y60VSS_X60Y70VSS X60Y65VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X60Y80VDD X60Y70VDD X60Y75VDD 25mOhm
L_X60Y70VDD_X60Y80VDD X60Y75VDD X60Y80VDD 2.91e-06nH
R_X60Y70VSS_X60Y80VSS X60Y70VSS X60Y75VSS 25mOhm
L_X60Y70VSS_X60Y80VSS X60Y75VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X60Y90VDD X60Y80VDD X60Y85VDD 25mOhm
L_X60Y80VDD_X60Y90VDD X60Y85VDD X60Y90VDD 2.91e-06nH
R_X60Y80VSS_X60Y90VSS X60Y80VSS X60Y85VSS 25mOhm
L_X60Y80VSS_X60Y90VSS X60Y85VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X60Y100VDD X60Y90VDD X60Y95VDD 25mOhm
L_X60Y90VDD_X60Y100VDD X60Y95VDD X60Y100VDD 2.91e-06nH
R_X60Y90VSS_X60Y100VSS X60Y90VSS X60Y95VSS 25mOhm
L_X60Y90VSS_X60Y100VSS X60Y95VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X60Y110VDD X60Y100VDD X60Y105VDD 25mOhm
L_X60Y100VDD_X60Y110VDD X60Y105VDD X60Y110VDD 2.91e-06nH
R_X60Y100VSS_X60Y110VSS X60Y100VSS X60Y105VSS 25mOhm
L_X60Y100VSS_X60Y110VSS X60Y105VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X60Y120VDD X60Y110VDD X60Y115VDD 25mOhm
L_X60Y110VDD_X60Y120VDD X60Y115VDD X60Y120VDD 2.91e-06nH
R_X60Y110VSS_X60Y120VSS X60Y110VSS X60Y115VSS 25mOhm
L_X60Y110VSS_X60Y120VSS X60Y115VSS X60Y120VSS 2.91e-06nH
R_X70Y10VDD_X70Y20VDD X70Y10VDD X70Y15VDD 25mOhm
L_X70Y10VDD_X70Y20VDD X70Y15VDD X70Y20VDD 2.91e-06nH
R_X70Y10VSS_X70Y20VSS X70Y10VSS X70Y15VSS 25mOhm
L_X70Y10VSS_X70Y20VSS X70Y15VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X70Y30VDD X70Y20VDD X70Y25VDD 25mOhm
L_X70Y20VDD_X70Y30VDD X70Y25VDD X70Y30VDD 2.91e-06nH
R_X70Y20VSS_X70Y30VSS X70Y20VSS X70Y25VSS 25mOhm
L_X70Y20VSS_X70Y30VSS X70Y25VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X70Y40VDD X70Y30VDD X70Y35VDD 25mOhm
L_X70Y30VDD_X70Y40VDD X70Y35VDD X70Y40VDD 2.91e-06nH
R_X70Y30VSS_X70Y40VSS X70Y30VSS X70Y35VSS 25mOhm
L_X70Y30VSS_X70Y40VSS X70Y35VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X70Y50VDD X70Y40VDD X70Y45VDD 25mOhm
L_X70Y40VDD_X70Y50VDD X70Y45VDD X70Y50VDD 2.91e-06nH
R_X70Y40VSS_X70Y50VSS X70Y40VSS X70Y45VSS 25mOhm
L_X70Y40VSS_X70Y50VSS X70Y45VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X70Y60VDD X70Y50VDD X70Y55VDD 25mOhm
L_X70Y50VDD_X70Y60VDD X70Y55VDD X70Y60VDD 2.91e-06nH
R_X70Y50VSS_X70Y60VSS X70Y50VSS X70Y55VSS 25mOhm
L_X70Y50VSS_X70Y60VSS X70Y55VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X70Y70VDD X70Y60VDD X70Y65VDD 25mOhm
L_X70Y60VDD_X70Y70VDD X70Y65VDD X70Y70VDD 2.91e-06nH
R_X70Y60VSS_X70Y70VSS X70Y60VSS X70Y65VSS 25mOhm
L_X70Y60VSS_X70Y70VSS X70Y65VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X70Y80VDD X70Y70VDD X70Y75VDD 25mOhm
L_X70Y70VDD_X70Y80VDD X70Y75VDD X70Y80VDD 2.91e-06nH
R_X70Y70VSS_X70Y80VSS X70Y70VSS X70Y75VSS 25mOhm
L_X70Y70VSS_X70Y80VSS X70Y75VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X70Y90VDD X70Y80VDD X70Y85VDD 25mOhm
L_X70Y80VDD_X70Y90VDD X70Y85VDD X70Y90VDD 2.91e-06nH
R_X70Y80VSS_X70Y90VSS X70Y80VSS X70Y85VSS 25mOhm
L_X70Y80VSS_X70Y90VSS X70Y85VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X70Y100VDD X70Y90VDD X70Y95VDD 25mOhm
L_X70Y90VDD_X70Y100VDD X70Y95VDD X70Y100VDD 2.91e-06nH
R_X70Y90VSS_X70Y100VSS X70Y90VSS X70Y95VSS 25mOhm
L_X70Y90VSS_X70Y100VSS X70Y95VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X70Y110VDD X70Y100VDD X70Y105VDD 25mOhm
L_X70Y100VDD_X70Y110VDD X70Y105VDD X70Y110VDD 2.91e-06nH
R_X70Y100VSS_X70Y110VSS X70Y100VSS X70Y105VSS 25mOhm
L_X70Y100VSS_X70Y110VSS X70Y105VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X70Y120VDD X70Y110VDD X70Y115VDD 25mOhm
L_X70Y110VDD_X70Y120VDD X70Y115VDD X70Y120VDD 2.91e-06nH
R_X70Y110VSS_X70Y120VSS X70Y110VSS X70Y115VSS 25mOhm
L_X70Y110VSS_X70Y120VSS X70Y115VSS X70Y120VSS 2.91e-06nH
R_X80Y10VDD_X80Y20VDD X80Y10VDD X80Y15VDD 25mOhm
L_X80Y10VDD_X80Y20VDD X80Y15VDD X80Y20VDD 2.91e-06nH
R_X80Y10VSS_X80Y20VSS X80Y10VSS X80Y15VSS 25mOhm
L_X80Y10VSS_X80Y20VSS X80Y15VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X80Y30VDD X80Y20VDD X80Y25VDD 25mOhm
L_X80Y20VDD_X80Y30VDD X80Y25VDD X80Y30VDD 2.91e-06nH
R_X80Y20VSS_X80Y30VSS X80Y20VSS X80Y25VSS 25mOhm
L_X80Y20VSS_X80Y30VSS X80Y25VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X80Y40VDD X80Y30VDD X80Y35VDD 25mOhm
L_X80Y30VDD_X80Y40VDD X80Y35VDD X80Y40VDD 2.91e-06nH
R_X80Y30VSS_X80Y40VSS X80Y30VSS X80Y35VSS 25mOhm
L_X80Y30VSS_X80Y40VSS X80Y35VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X80Y50VDD X80Y40VDD X80Y45VDD 25mOhm
L_X80Y40VDD_X80Y50VDD X80Y45VDD X80Y50VDD 2.91e-06nH
R_X80Y40VSS_X80Y50VSS X80Y40VSS X80Y45VSS 25mOhm
L_X80Y40VSS_X80Y50VSS X80Y45VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X80Y60VDD X80Y50VDD X80Y55VDD 25mOhm
L_X80Y50VDD_X80Y60VDD X80Y55VDD X80Y60VDD 2.91e-06nH
R_X80Y50VSS_X80Y60VSS X80Y50VSS X80Y55VSS 25mOhm
L_X80Y50VSS_X80Y60VSS X80Y55VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X80Y70VDD X80Y60VDD X80Y65VDD 25mOhm
L_X80Y60VDD_X80Y70VDD X80Y65VDD X80Y70VDD 2.91e-06nH
R_X80Y60VSS_X80Y70VSS X80Y60VSS X80Y65VSS 25mOhm
L_X80Y60VSS_X80Y70VSS X80Y65VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X80Y80VDD X80Y70VDD X80Y75VDD 25mOhm
L_X80Y70VDD_X80Y80VDD X80Y75VDD X80Y80VDD 2.91e-06nH
R_X80Y70VSS_X80Y80VSS X80Y70VSS X80Y75VSS 25mOhm
L_X80Y70VSS_X80Y80VSS X80Y75VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X80Y90VDD X80Y80VDD X80Y85VDD 25mOhm
L_X80Y80VDD_X80Y90VDD X80Y85VDD X80Y90VDD 2.91e-06nH
R_X80Y80VSS_X80Y90VSS X80Y80VSS X80Y85VSS 25mOhm
L_X80Y80VSS_X80Y90VSS X80Y85VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X80Y100VDD X80Y90VDD X80Y95VDD 25mOhm
L_X80Y90VDD_X80Y100VDD X80Y95VDD X80Y100VDD 2.91e-06nH
R_X80Y90VSS_X80Y100VSS X80Y90VSS X80Y95VSS 25mOhm
L_X80Y90VSS_X80Y100VSS X80Y95VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X80Y110VDD X80Y100VDD X80Y105VDD 25mOhm
L_X80Y100VDD_X80Y110VDD X80Y105VDD X80Y110VDD 2.91e-06nH
R_X80Y100VSS_X80Y110VSS X80Y100VSS X80Y105VSS 25mOhm
L_X80Y100VSS_X80Y110VSS X80Y105VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X80Y120VDD X80Y110VDD X80Y115VDD 25mOhm
L_X80Y110VDD_X80Y120VDD X80Y115VDD X80Y120VDD 2.91e-06nH
R_X80Y110VSS_X80Y120VSS X80Y110VSS X80Y115VSS 25mOhm
L_X80Y110VSS_X80Y120VSS X80Y115VSS X80Y120VSS 2.91e-06nH
R_X90Y10VDD_X90Y20VDD X90Y10VDD X90Y15VDD 25mOhm
L_X90Y10VDD_X90Y20VDD X90Y15VDD X90Y20VDD 2.91e-06nH
R_X90Y10VSS_X90Y20VSS X90Y10VSS X90Y15VSS 25mOhm
L_X90Y10VSS_X90Y20VSS X90Y15VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X90Y30VDD X90Y20VDD X90Y25VDD 25mOhm
L_X90Y20VDD_X90Y30VDD X90Y25VDD X90Y30VDD 2.91e-06nH
R_X90Y20VSS_X90Y30VSS X90Y20VSS X90Y25VSS 25mOhm
L_X90Y20VSS_X90Y30VSS X90Y25VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X90Y40VDD X90Y30VDD X90Y35VDD 25mOhm
L_X90Y30VDD_X90Y40VDD X90Y35VDD X90Y40VDD 2.91e-06nH
R_X90Y30VSS_X90Y40VSS X90Y30VSS X90Y35VSS 25mOhm
L_X90Y30VSS_X90Y40VSS X90Y35VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X90Y50VDD X90Y40VDD X90Y45VDD 25mOhm
L_X90Y40VDD_X90Y50VDD X90Y45VDD X90Y50VDD 2.91e-06nH
R_X90Y40VSS_X90Y50VSS X90Y40VSS X90Y45VSS 25mOhm
L_X90Y40VSS_X90Y50VSS X90Y45VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X90Y60VDD X90Y50VDD X90Y55VDD 25mOhm
L_X90Y50VDD_X90Y60VDD X90Y55VDD X90Y60VDD 2.91e-06nH
R_X90Y50VSS_X90Y60VSS X90Y50VSS X90Y55VSS 25mOhm
L_X90Y50VSS_X90Y60VSS X90Y55VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X90Y70VDD X90Y60VDD X90Y65VDD 25mOhm
L_X90Y60VDD_X90Y70VDD X90Y65VDD X90Y70VDD 2.91e-06nH
R_X90Y60VSS_X90Y70VSS X90Y60VSS X90Y65VSS 25mOhm
L_X90Y60VSS_X90Y70VSS X90Y65VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X90Y80VDD X90Y70VDD X90Y75VDD 25mOhm
L_X90Y70VDD_X90Y80VDD X90Y75VDD X90Y80VDD 2.91e-06nH
R_X90Y70VSS_X90Y80VSS X90Y70VSS X90Y75VSS 25mOhm
L_X90Y70VSS_X90Y80VSS X90Y75VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X90Y90VDD X90Y80VDD X90Y85VDD 25mOhm
L_X90Y80VDD_X90Y90VDD X90Y85VDD X90Y90VDD 2.91e-06nH
R_X90Y80VSS_X90Y90VSS X90Y80VSS X90Y85VSS 25mOhm
L_X90Y80VSS_X90Y90VSS X90Y85VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X90Y100VDD X90Y90VDD X90Y95VDD 25mOhm
L_X90Y90VDD_X90Y100VDD X90Y95VDD X90Y100VDD 2.91e-06nH
R_X90Y90VSS_X90Y100VSS X90Y90VSS X90Y95VSS 25mOhm
L_X90Y90VSS_X90Y100VSS X90Y95VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X90Y110VDD X90Y100VDD X90Y105VDD 25mOhm
L_X90Y100VDD_X90Y110VDD X90Y105VDD X90Y110VDD 2.91e-06nH
R_X90Y100VSS_X90Y110VSS X90Y100VSS X90Y105VSS 25mOhm
L_X90Y100VSS_X90Y110VSS X90Y105VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X90Y120VDD X90Y110VDD X90Y115VDD 25mOhm
L_X90Y110VDD_X90Y120VDD X90Y115VDD X90Y120VDD 2.91e-06nH
R_X90Y110VSS_X90Y120VSS X90Y110VSS X90Y115VSS 25mOhm
L_X90Y110VSS_X90Y120VSS X90Y115VSS X90Y120VSS 2.91e-06nH
R_X100Y10VDD_X100Y20VDD X100Y10VDD X100Y15VDD 25mOhm
L_X100Y10VDD_X100Y20VDD X100Y15VDD X100Y20VDD 2.91e-06nH
R_X100Y10VSS_X100Y20VSS X100Y10VSS X100Y15VSS 25mOhm
L_X100Y10VSS_X100Y20VSS X100Y15VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X100Y30VDD X100Y20VDD X100Y25VDD 25mOhm
L_X100Y20VDD_X100Y30VDD X100Y25VDD X100Y30VDD 2.91e-06nH
R_X100Y20VSS_X100Y30VSS X100Y20VSS X100Y25VSS 25mOhm
L_X100Y20VSS_X100Y30VSS X100Y25VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X100Y40VDD X100Y30VDD X100Y35VDD 25mOhm
L_X100Y30VDD_X100Y40VDD X100Y35VDD X100Y40VDD 2.91e-06nH
R_X100Y30VSS_X100Y40VSS X100Y30VSS X100Y35VSS 25mOhm
L_X100Y30VSS_X100Y40VSS X100Y35VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X100Y50VDD X100Y40VDD X100Y45VDD 25mOhm
L_X100Y40VDD_X100Y50VDD X100Y45VDD X100Y50VDD 2.91e-06nH
R_X100Y40VSS_X100Y50VSS X100Y40VSS X100Y45VSS 25mOhm
L_X100Y40VSS_X100Y50VSS X100Y45VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X100Y60VDD X100Y50VDD X100Y55VDD 25mOhm
L_X100Y50VDD_X100Y60VDD X100Y55VDD X100Y60VDD 2.91e-06nH
R_X100Y50VSS_X100Y60VSS X100Y50VSS X100Y55VSS 25mOhm
L_X100Y50VSS_X100Y60VSS X100Y55VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X100Y70VDD X100Y60VDD X100Y65VDD 25mOhm
L_X100Y60VDD_X100Y70VDD X100Y65VDD X100Y70VDD 2.91e-06nH
R_X100Y60VSS_X100Y70VSS X100Y60VSS X100Y65VSS 25mOhm
L_X100Y60VSS_X100Y70VSS X100Y65VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X100Y80VDD X100Y70VDD X100Y75VDD 25mOhm
L_X100Y70VDD_X100Y80VDD X100Y75VDD X100Y80VDD 2.91e-06nH
R_X100Y70VSS_X100Y80VSS X100Y70VSS X100Y75VSS 25mOhm
L_X100Y70VSS_X100Y80VSS X100Y75VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X100Y90VDD X100Y80VDD X100Y85VDD 25mOhm
L_X100Y80VDD_X100Y90VDD X100Y85VDD X100Y90VDD 2.91e-06nH
R_X100Y80VSS_X100Y90VSS X100Y80VSS X100Y85VSS 25mOhm
L_X100Y80VSS_X100Y90VSS X100Y85VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X100Y100VDD X100Y90VDD X100Y95VDD 25mOhm
L_X100Y90VDD_X100Y100VDD X100Y95VDD X100Y100VDD 2.91e-06nH
R_X100Y90VSS_X100Y100VSS X100Y90VSS X100Y95VSS 25mOhm
L_X100Y90VSS_X100Y100VSS X100Y95VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X100Y110VDD X100Y100VDD X100Y105VDD 25mOhm
L_X100Y100VDD_X100Y110VDD X100Y105VDD X100Y110VDD 2.91e-06nH
R_X100Y100VSS_X100Y110VSS X100Y100VSS X100Y105VSS 25mOhm
L_X100Y100VSS_X100Y110VSS X100Y105VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X100Y120VDD X100Y110VDD X100Y115VDD 25mOhm
L_X100Y110VDD_X100Y120VDD X100Y115VDD X100Y120VDD 2.91e-06nH
R_X100Y110VSS_X100Y120VSS X100Y110VSS X100Y115VSS 25mOhm
L_X100Y110VSS_X100Y120VSS X100Y115VSS X100Y120VSS 2.91e-06nH
R_X110Y10VDD_X110Y20VDD X110Y10VDD X110Y15VDD 25mOhm
L_X110Y10VDD_X110Y20VDD X110Y15VDD X110Y20VDD 2.91e-06nH
R_X110Y10VSS_X110Y20VSS X110Y10VSS X110Y15VSS 25mOhm
L_X110Y10VSS_X110Y20VSS X110Y15VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X110Y30VDD X110Y20VDD X110Y25VDD 25mOhm
L_X110Y20VDD_X110Y30VDD X110Y25VDD X110Y30VDD 2.91e-06nH
R_X110Y20VSS_X110Y30VSS X110Y20VSS X110Y25VSS 25mOhm
L_X110Y20VSS_X110Y30VSS X110Y25VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X110Y40VDD X110Y30VDD X110Y35VDD 25mOhm
L_X110Y30VDD_X110Y40VDD X110Y35VDD X110Y40VDD 2.91e-06nH
R_X110Y30VSS_X110Y40VSS X110Y30VSS X110Y35VSS 25mOhm
L_X110Y30VSS_X110Y40VSS X110Y35VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X110Y50VDD X110Y40VDD X110Y45VDD 25mOhm
L_X110Y40VDD_X110Y50VDD X110Y45VDD X110Y50VDD 2.91e-06nH
R_X110Y40VSS_X110Y50VSS X110Y40VSS X110Y45VSS 25mOhm
L_X110Y40VSS_X110Y50VSS X110Y45VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X110Y60VDD X110Y50VDD X110Y55VDD 25mOhm
L_X110Y50VDD_X110Y60VDD X110Y55VDD X110Y60VDD 2.91e-06nH
R_X110Y50VSS_X110Y60VSS X110Y50VSS X110Y55VSS 25mOhm
L_X110Y50VSS_X110Y60VSS X110Y55VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X110Y70VDD X110Y60VDD X110Y65VDD 25mOhm
L_X110Y60VDD_X110Y70VDD X110Y65VDD X110Y70VDD 2.91e-06nH
R_X110Y60VSS_X110Y70VSS X110Y60VSS X110Y65VSS 25mOhm
L_X110Y60VSS_X110Y70VSS X110Y65VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X110Y80VDD X110Y70VDD X110Y75VDD 25mOhm
L_X110Y70VDD_X110Y80VDD X110Y75VDD X110Y80VDD 2.91e-06nH
R_X110Y70VSS_X110Y80VSS X110Y70VSS X110Y75VSS 25mOhm
L_X110Y70VSS_X110Y80VSS X110Y75VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X110Y90VDD X110Y80VDD X110Y85VDD 25mOhm
L_X110Y80VDD_X110Y90VDD X110Y85VDD X110Y90VDD 2.91e-06nH
R_X110Y80VSS_X110Y90VSS X110Y80VSS X110Y85VSS 25mOhm
L_X110Y80VSS_X110Y90VSS X110Y85VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X110Y100VDD X110Y90VDD X110Y95VDD 25mOhm
L_X110Y90VDD_X110Y100VDD X110Y95VDD X110Y100VDD 2.91e-06nH
R_X110Y90VSS_X110Y100VSS X110Y90VSS X110Y95VSS 25mOhm
L_X110Y90VSS_X110Y100VSS X110Y95VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X110Y110VDD X110Y100VDD X110Y105VDD 25mOhm
L_X110Y100VDD_X110Y110VDD X110Y105VDD X110Y110VDD 2.91e-06nH
R_X110Y100VSS_X110Y110VSS X110Y100VSS X110Y105VSS 25mOhm
L_X110Y100VSS_X110Y110VSS X110Y105VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X110Y120VDD X110Y110VDD X110Y115VDD 25mOhm
L_X110Y110VDD_X110Y120VDD X110Y115VDD X110Y120VDD 2.91e-06nH
R_X110Y110VSS_X110Y120VSS X110Y110VSS X110Y115VSS 25mOhm
L_X110Y110VSS_X110Y120VSS X110Y115VSS X110Y120VSS 2.91e-06nH
R_X120Y10VDD_X120Y20VDD X120Y10VDD X120Y15VDD 25mOhm
L_X120Y10VDD_X120Y20VDD X120Y15VDD X120Y20VDD 2.91e-06nH
R_X120Y10VSS_X120Y20VSS X120Y10VSS X120Y15VSS 25mOhm
L_X120Y10VSS_X120Y20VSS X120Y15VSS X120Y20VSS 2.91e-06nH
R_X120Y20VDD_X120Y30VDD X120Y20VDD X120Y25VDD 25mOhm
L_X120Y20VDD_X120Y30VDD X120Y25VDD X120Y30VDD 2.91e-06nH
R_X120Y20VSS_X120Y30VSS X120Y20VSS X120Y25VSS 25mOhm
L_X120Y20VSS_X120Y30VSS X120Y25VSS X120Y30VSS 2.91e-06nH
R_X120Y30VDD_X120Y40VDD X120Y30VDD X120Y35VDD 25mOhm
L_X120Y30VDD_X120Y40VDD X120Y35VDD X120Y40VDD 2.91e-06nH
R_X120Y30VSS_X120Y40VSS X120Y30VSS X120Y35VSS 25mOhm
L_X120Y30VSS_X120Y40VSS X120Y35VSS X120Y40VSS 2.91e-06nH
R_X120Y40VDD_X120Y50VDD X120Y40VDD X120Y45VDD 25mOhm
L_X120Y40VDD_X120Y50VDD X120Y45VDD X120Y50VDD 2.91e-06nH
R_X120Y40VSS_X120Y50VSS X120Y40VSS X120Y45VSS 25mOhm
L_X120Y40VSS_X120Y50VSS X120Y45VSS X120Y50VSS 2.91e-06nH
R_X120Y50VDD_X120Y60VDD X120Y50VDD X120Y55VDD 25mOhm
L_X120Y50VDD_X120Y60VDD X120Y55VDD X120Y60VDD 2.91e-06nH
R_X120Y50VSS_X120Y60VSS X120Y50VSS X120Y55VSS 25mOhm
L_X120Y50VSS_X120Y60VSS X120Y55VSS X120Y60VSS 2.91e-06nH
R_X120Y60VDD_X120Y70VDD X120Y60VDD X120Y65VDD 25mOhm
L_X120Y60VDD_X120Y70VDD X120Y65VDD X120Y70VDD 2.91e-06nH
R_X120Y60VSS_X120Y70VSS X120Y60VSS X120Y65VSS 25mOhm
L_X120Y60VSS_X120Y70VSS X120Y65VSS X120Y70VSS 2.91e-06nH
R_X120Y70VDD_X120Y80VDD X120Y70VDD X120Y75VDD 25mOhm
L_X120Y70VDD_X120Y80VDD X120Y75VDD X120Y80VDD 2.91e-06nH
R_X120Y70VSS_X120Y80VSS X120Y70VSS X120Y75VSS 25mOhm
L_X120Y70VSS_X120Y80VSS X120Y75VSS X120Y80VSS 2.91e-06nH
R_X120Y80VDD_X120Y90VDD X120Y80VDD X120Y85VDD 25mOhm
L_X120Y80VDD_X120Y90VDD X120Y85VDD X120Y90VDD 2.91e-06nH
R_X120Y80VSS_X120Y90VSS X120Y80VSS X120Y85VSS 25mOhm
L_X120Y80VSS_X120Y90VSS X120Y85VSS X120Y90VSS 2.91e-06nH
R_X120Y90VDD_X120Y100VDD X120Y90VDD X120Y95VDD 25mOhm
L_X120Y90VDD_X120Y100VDD X120Y95VDD X120Y100VDD 2.91e-06nH
R_X120Y90VSS_X120Y100VSS X120Y90VSS X120Y95VSS 25mOhm
L_X120Y90VSS_X120Y100VSS X120Y95VSS X120Y100VSS 2.91e-06nH
R_X120Y100VDD_X120Y110VDD X120Y100VDD X120Y105VDD 25mOhm
L_X120Y100VDD_X120Y110VDD X120Y105VDD X120Y110VDD 2.91e-06nH
R_X120Y100VSS_X120Y110VSS X120Y100VSS X120Y105VSS 25mOhm
L_X120Y100VSS_X120Y110VSS X120Y105VSS X120Y110VSS 2.91e-06nH
R_X120Y110VDD_X120Y120VDD X120Y110VDD X120Y115VDD 25mOhm
L_X120Y110VDD_X120Y120VDD X120Y115VDD X120Y120VDD 2.91e-06nH
R_X120Y110VSS_X120Y120VSS X120Y110VSS X120Y115VSS 25mOhm
L_X120Y110VSS_X120Y120VSS X120Y115VSS X120Y120VSS 2.91e-06nH
C_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VSS 10nF
C_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VSS 10nF
C_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VSS 10nF
C_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VSS 10nF
C_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VSS 10nF
C_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VSS 10nF
C_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VSS 10nF
C_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VSS 10nF
C_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VSS 10nF
C_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VSS 10nF
C_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VSS 10nF
C_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VSS 10nF
C_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VSS 10nF
C_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VSS 10nF
C_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VSS 10nF
C_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VSS 10nF
C_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VSS 10nF
C_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VSS 10nF
C_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VSS 10nF
C_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VSS 10nF
C_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VSS 10nF
C_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VSS 10nF
C_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VSS 10nF
C_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VSS 10nF
C_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VSS 10nF
C_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VSS 10nF
C_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VSS 10nF
C_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VSS 10nF
C_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VSS 10nF
C_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VSS 10nF
C_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VSS 10nF
C_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VSS 10nF
C_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VSS 10nF
C_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VSS 10nF
C_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VSS 10nF
C_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VSS 10nF
C_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VSS 10nF
C_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VSS 10nF
C_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VSS 10nF
C_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VSS 10nF
C_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VSS 10nF
C_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VSS 10nF
C_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VSS 10nF
C_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VSS 10nF
C_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VSS 10nF
C_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VSS 10nF
C_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VSS 10nF
C_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VSS 10nF
C_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VSS 10nF
C_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VSS 10nF
C_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VSS 10nF
C_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VSS 10nF
C_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VSS 10nF
C_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VSS 10nF
C_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VSS 10nF
C_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VSS 10nF
C_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VSS 10nF
C_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VSS 10nF
C_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VSS 10nF
C_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VSS 10nF
C_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VSS 10nF
C_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VSS 10nF
C_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VSS 10nF
C_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VSS 10nF
C_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VSS 10nF
C_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VSS 10nF
C_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VSS 10nF
C_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VSS 10nF
C_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VSS 10nF
C_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VSS 10nF
C_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VSS 10nF
C_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VSS 10nF
C_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VSS 10nF
C_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VSS 10nF
C_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VSS 10nF
C_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VSS 10nF
C_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VSS 10nF
C_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VSS 10nF
C_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VSS 10nF
C_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VSS 10nF
C_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VSS 10nF
C_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VSS 10nF
C_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VSS 10nF
C_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VSS 10nF
C_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VSS 10nF
C_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VSS 10nF
C_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VSS 10nF
C_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VSS 10nF
C_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VSS 10nF
C_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VSS 10nF
C_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VSS 10nF
C_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VSS 10nF
C_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VSS 10nF
C_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VSS 10nF
C_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VSS 10nF
C_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VSS 10nF
C_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VSS 10nF
C_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VSS 10nF
C_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VSS 10nF
C_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VSS 10nF
C_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VSS 10nF
C_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VSS 10nF
C_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VSS 10nF
C_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VSS 10nF
C_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VSS 10nF
C_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VSS 10nF
C_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VSS 10nF
C_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VSS 10nF
C_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VSS 10nF
C_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VSS 10nF
C_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VSS 10nF
C_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VSS 10nF
C_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VSS 10nF
C_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VSS 10nF
C_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VSS 10nF
C_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VSS 10nF
C_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VSS 10nF
C_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VSS 10nF
C_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VSS 10nF
C_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VSS 10nF
C_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VSS 10nF
C_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VSS 10nF
C_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VSS 10nF
C_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VSS 10nF
C_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VSS 10nF
C_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VSS 10nF
C_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VSS 10nF
C_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VSS 10nF
C_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VSS 10nF
C_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VSS 10nF
C_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VSS 10nF
C_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VSS 10nF
C_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VSS 10nF
C_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VSS 10nF
C_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VSS 10nF
C_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VSS 10nF
C_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VSS 10nF
C_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VSS 10nF
C_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VSS 10nF
C_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VSS 10nF
C_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VSS 10nF
C_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VSS 10nF
C_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VSS 10nF
C_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VSS 10nF
I_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VDDDM 1 AC=0.006944444444444444
V_X120Y120VDD_X120Y120VSS X120Y120VDDDM X120Y120VSS 0
I_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VDDDM 1 AC=0.006944444444444444
V_X120Y10VDD_X120Y10VSS X120Y10VDDDM X120Y10VSS 0
I_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VDDDM 1 AC=0.006944444444444444
V_X120Y20VDD_X120Y20VSS X120Y20VDDDM X120Y20VSS 0
I_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VDDDM 1 AC=0.006944444444444444
V_X120Y30VDD_X120Y30VSS X120Y30VDDDM X120Y30VSS 0
I_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VDDDM 1 AC=0.006944444444444444
V_X120Y40VDD_X120Y40VSS X120Y40VDDDM X120Y40VSS 0
I_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VDDDM 1 AC=0.006944444444444444
V_X120Y50VDD_X120Y50VSS X120Y50VDDDM X120Y50VSS 0
I_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VDDDM 1 AC=0.006944444444444444
V_X120Y60VDD_X120Y60VSS X120Y60VDDDM X120Y60VSS 0
I_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VDDDM 1 AC=0.006944444444444444
V_X120Y70VDD_X120Y70VSS X120Y70VDDDM X120Y70VSS 0
I_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VDDDM 1 AC=0.006944444444444444
V_X120Y80VDD_X120Y80VSS X120Y80VDDDM X120Y80VSS 0
I_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VDDDM 1 AC=0.006944444444444444
V_X120Y90VDD_X120Y90VSS X120Y90VDDDM X120Y90VSS 0
I_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VDDDM 1 AC=0.006944444444444444
V_X120Y100VDD_X120Y100VSS X120Y100VDDDM X120Y100VSS 0
I_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VDDDM 1 AC=0.006944444444444444
V_X120Y110VDD_X120Y110VSS X120Y110VDDDM X120Y110VSS 0
I_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VDDDM 1 AC=0.006944444444444444
V_X10Y120VDD_X10Y120VSS X10Y120VDDDM X10Y120VSS 0
I_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VDDDM 1 AC=0.006944444444444444
V_X10Y10VDD_X10Y10VSS X10Y10VDDDM X10Y10VSS 0
I_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VDDDM 1 AC=0.006944444444444444
V_X10Y20VDD_X10Y20VSS X10Y20VDDDM X10Y20VSS 0
I_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VDDDM 1 AC=0.006944444444444444
V_X10Y30VDD_X10Y30VSS X10Y30VDDDM X10Y30VSS 0
I_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VDDDM 1 AC=0.006944444444444444
V_X10Y40VDD_X10Y40VSS X10Y40VDDDM X10Y40VSS 0
I_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VDDDM 1 AC=0.006944444444444444
V_X10Y50VDD_X10Y50VSS X10Y50VDDDM X10Y50VSS 0
I_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VDDDM 1 AC=0.006944444444444444
V_X10Y60VDD_X10Y60VSS X10Y60VDDDM X10Y60VSS 0
I_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VDDDM 1 AC=0.006944444444444444
V_X10Y70VDD_X10Y70VSS X10Y70VDDDM X10Y70VSS 0
I_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VDDDM 1 AC=0.006944444444444444
V_X10Y80VDD_X10Y80VSS X10Y80VDDDM X10Y80VSS 0
I_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VDDDM 1 AC=0.006944444444444444
V_X10Y90VDD_X10Y90VSS X10Y90VDDDM X10Y90VSS 0
I_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VDDDM 1 AC=0.006944444444444444
V_X10Y100VDD_X10Y100VSS X10Y100VDDDM X10Y100VSS 0
I_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VDDDM 1 AC=0.006944444444444444
V_X10Y110VDD_X10Y110VSS X10Y110VDDDM X10Y110VSS 0
I_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VDDDM 1 AC=0.006944444444444444
V_X20Y120VDD_X20Y120VSS X20Y120VDDDM X20Y120VSS 0
I_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VDDDM 1 AC=0.006944444444444444
V_X20Y10VDD_X20Y10VSS X20Y10VDDDM X20Y10VSS 0
I_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VDDDM 1 AC=0.006944444444444444
V_X20Y20VDD_X20Y20VSS X20Y20VDDDM X20Y20VSS 0
I_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VDDDM 1 AC=0.006944444444444444
V_X20Y30VDD_X20Y30VSS X20Y30VDDDM X20Y30VSS 0
I_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VDDDM 1 AC=0.006944444444444444
V_X20Y40VDD_X20Y40VSS X20Y40VDDDM X20Y40VSS 0
I_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VDDDM 1 AC=0.006944444444444444
V_X20Y50VDD_X20Y50VSS X20Y50VDDDM X20Y50VSS 0
I_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VDDDM 1 AC=0.006944444444444444
V_X20Y60VDD_X20Y60VSS X20Y60VDDDM X20Y60VSS 0
I_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VDDDM 1 AC=0.006944444444444444
V_X20Y70VDD_X20Y70VSS X20Y70VDDDM X20Y70VSS 0
I_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VDDDM 1 AC=0.006944444444444444
V_X20Y80VDD_X20Y80VSS X20Y80VDDDM X20Y80VSS 0
I_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VDDDM 1 AC=0.006944444444444444
V_X20Y90VDD_X20Y90VSS X20Y90VDDDM X20Y90VSS 0
I_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VDDDM 1 AC=0.006944444444444444
V_X20Y100VDD_X20Y100VSS X20Y100VDDDM X20Y100VSS 0
I_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VDDDM 1 AC=0.006944444444444444
V_X20Y110VDD_X20Y110VSS X20Y110VDDDM X20Y110VSS 0
I_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VDDDM 1 AC=0.006944444444444444
V_X30Y120VDD_X30Y120VSS X30Y120VDDDM X30Y120VSS 0
I_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VDDDM 1 AC=0.006944444444444444
V_X30Y10VDD_X30Y10VSS X30Y10VDDDM X30Y10VSS 0
I_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VDDDM 1 AC=0.006944444444444444
V_X30Y20VDD_X30Y20VSS X30Y20VDDDM X30Y20VSS 0
I_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VDDDM 1 AC=0.006944444444444444
V_X30Y30VDD_X30Y30VSS X30Y30VDDDM X30Y30VSS 0
I_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VDDDM 1 AC=0.006944444444444444
V_X30Y40VDD_X30Y40VSS X30Y40VDDDM X30Y40VSS 0
I_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VDDDM 1 AC=0.006944444444444444
V_X30Y50VDD_X30Y50VSS X30Y50VDDDM X30Y50VSS 0
I_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VDDDM 1 AC=0.006944444444444444
V_X30Y60VDD_X30Y60VSS X30Y60VDDDM X30Y60VSS 0
I_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VDDDM 1 AC=0.006944444444444444
V_X30Y70VDD_X30Y70VSS X30Y70VDDDM X30Y70VSS 0
I_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VDDDM 1 AC=0.006944444444444444
V_X30Y80VDD_X30Y80VSS X30Y80VDDDM X30Y80VSS 0
I_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VDDDM 1 AC=0.006944444444444444
V_X30Y90VDD_X30Y90VSS X30Y90VDDDM X30Y90VSS 0
I_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VDDDM 1 AC=0.006944444444444444
V_X30Y100VDD_X30Y100VSS X30Y100VDDDM X30Y100VSS 0
I_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VDDDM 1 AC=0.006944444444444444
V_X30Y110VDD_X30Y110VSS X30Y110VDDDM X30Y110VSS 0
I_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VDDDM 1 AC=0.006944444444444444
V_X40Y120VDD_X40Y120VSS X40Y120VDDDM X40Y120VSS 0
I_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VDDDM 1 AC=0.006944444444444444
V_X40Y10VDD_X40Y10VSS X40Y10VDDDM X40Y10VSS 0
I_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VDDDM 1 AC=0.006944444444444444
V_X40Y20VDD_X40Y20VSS X40Y20VDDDM X40Y20VSS 0
I_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VDDDM 1 AC=0.006944444444444444
V_X40Y30VDD_X40Y30VSS X40Y30VDDDM X40Y30VSS 0
I_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VDDDM 1 AC=0.006944444444444444
V_X40Y40VDD_X40Y40VSS X40Y40VDDDM X40Y40VSS 0
I_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VDDDM 1 AC=0.006944444444444444
V_X40Y50VDD_X40Y50VSS X40Y50VDDDM X40Y50VSS 0
I_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VDDDM 1 AC=0.006944444444444444
V_X40Y60VDD_X40Y60VSS X40Y60VDDDM X40Y60VSS 0
I_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VDDDM 1 AC=0.006944444444444444
V_X40Y70VDD_X40Y70VSS X40Y70VDDDM X40Y70VSS 0
I_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VDDDM 1 AC=0.006944444444444444
V_X40Y80VDD_X40Y80VSS X40Y80VDDDM X40Y80VSS 0
I_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VDDDM 1 AC=0.006944444444444444
V_X40Y90VDD_X40Y90VSS X40Y90VDDDM X40Y90VSS 0
I_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VDDDM 1 AC=0.006944444444444444
V_X40Y100VDD_X40Y100VSS X40Y100VDDDM X40Y100VSS 0
I_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VDDDM 1 AC=0.006944444444444444
V_X40Y110VDD_X40Y110VSS X40Y110VDDDM X40Y110VSS 0
I_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VDDDM 1 AC=0.006944444444444444
V_X50Y120VDD_X50Y120VSS X50Y120VDDDM X50Y120VSS 0
I_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VDDDM 1 AC=0.006944444444444444
V_X50Y10VDD_X50Y10VSS X50Y10VDDDM X50Y10VSS 0
I_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VDDDM 1 AC=0.006944444444444444
V_X50Y20VDD_X50Y20VSS X50Y20VDDDM X50Y20VSS 0
I_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VDDDM 1 AC=0.006944444444444444
V_X50Y30VDD_X50Y30VSS X50Y30VDDDM X50Y30VSS 0
I_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VDDDM 1 AC=0.006944444444444444
V_X50Y40VDD_X50Y40VSS X50Y40VDDDM X50Y40VSS 0
I_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VDDDM 1 AC=0.006944444444444444
V_X50Y50VDD_X50Y50VSS X50Y50VDDDM X50Y50VSS 0
I_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VDDDM 1 AC=0.006944444444444444
V_X50Y60VDD_X50Y60VSS X50Y60VDDDM X50Y60VSS 0
I_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VDDDM 1 AC=0.006944444444444444
V_X50Y70VDD_X50Y70VSS X50Y70VDDDM X50Y70VSS 0
I_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VDDDM 1 AC=0.006944444444444444
V_X50Y80VDD_X50Y80VSS X50Y80VDDDM X50Y80VSS 0
I_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VDDDM 1 AC=0.006944444444444444
V_X50Y90VDD_X50Y90VSS X50Y90VDDDM X50Y90VSS 0
I_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VDDDM 1 AC=0.006944444444444444
V_X50Y100VDD_X50Y100VSS X50Y100VDDDM X50Y100VSS 0
I_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VDDDM 1 AC=0.006944444444444444
V_X50Y110VDD_X50Y110VSS X50Y110VDDDM X50Y110VSS 0
I_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VDDDM 1 AC=0.006944444444444444
V_X60Y120VDD_X60Y120VSS X60Y120VDDDM X60Y120VSS 0
I_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VDDDM 1 AC=0.006944444444444444
V_X60Y10VDD_X60Y10VSS X60Y10VDDDM X60Y10VSS 0
I_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VDDDM 1 AC=0.006944444444444444
V_X60Y20VDD_X60Y20VSS X60Y20VDDDM X60Y20VSS 0
I_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VDDDM 1 AC=0.006944444444444444
V_X60Y30VDD_X60Y30VSS X60Y30VDDDM X60Y30VSS 0
I_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VDDDM 1 AC=0.006944444444444444
V_X60Y40VDD_X60Y40VSS X60Y40VDDDM X60Y40VSS 0
I_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VDDDM 1 AC=0.006944444444444444
V_X60Y50VDD_X60Y50VSS X60Y50VDDDM X60Y50VSS 0
I_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VDDDM 1 AC=0.006944444444444444
V_X60Y60VDD_X60Y60VSS X60Y60VDDDM X60Y60VSS 0
I_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VDDDM 1 AC=0.006944444444444444
V_X60Y70VDD_X60Y70VSS X60Y70VDDDM X60Y70VSS 0
I_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VDDDM 1 AC=0.006944444444444444
V_X60Y80VDD_X60Y80VSS X60Y80VDDDM X60Y80VSS 0
I_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VDDDM 1 AC=0.006944444444444444
V_X60Y90VDD_X60Y90VSS X60Y90VDDDM X60Y90VSS 0
I_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VDDDM 1 AC=0.006944444444444444
V_X60Y100VDD_X60Y100VSS X60Y100VDDDM X60Y100VSS 0
I_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VDDDM 1 AC=0.006944444444444444
V_X60Y110VDD_X60Y110VSS X60Y110VDDDM X60Y110VSS 0
I_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VDDDM 1 AC=0.006944444444444444
V_X70Y120VDD_X70Y120VSS X70Y120VDDDM X70Y120VSS 0
I_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VDDDM 1 AC=0.006944444444444444
V_X70Y10VDD_X70Y10VSS X70Y10VDDDM X70Y10VSS 0
I_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VDDDM 1 AC=0.006944444444444444
V_X70Y20VDD_X70Y20VSS X70Y20VDDDM X70Y20VSS 0
I_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VDDDM 1 AC=0.006944444444444444
V_X70Y30VDD_X70Y30VSS X70Y30VDDDM X70Y30VSS 0
I_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VDDDM 1 AC=0.006944444444444444
V_X70Y40VDD_X70Y40VSS X70Y40VDDDM X70Y40VSS 0
I_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VDDDM 1 AC=0.006944444444444444
V_X70Y50VDD_X70Y50VSS X70Y50VDDDM X70Y50VSS 0
I_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VDDDM 1 AC=0.006944444444444444
V_X70Y60VDD_X70Y60VSS X70Y60VDDDM X70Y60VSS 0
I_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VDDDM 1 AC=0.006944444444444444
V_X70Y70VDD_X70Y70VSS X70Y70VDDDM X70Y70VSS 0
I_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VDDDM 1 AC=0.006944444444444444
V_X70Y80VDD_X70Y80VSS X70Y80VDDDM X70Y80VSS 0
I_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VDDDM 1 AC=0.006944444444444444
V_X70Y90VDD_X70Y90VSS X70Y90VDDDM X70Y90VSS 0
I_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VDDDM 1 AC=0.006944444444444444
V_X70Y100VDD_X70Y100VSS X70Y100VDDDM X70Y100VSS 0
I_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VDDDM 1 AC=0.006944444444444444
V_X70Y110VDD_X70Y110VSS X70Y110VDDDM X70Y110VSS 0
I_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VDDDM 1 AC=0.006944444444444444
V_X80Y120VDD_X80Y120VSS X80Y120VDDDM X80Y120VSS 0
I_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VDDDM 1 AC=0.006944444444444444
V_X80Y10VDD_X80Y10VSS X80Y10VDDDM X80Y10VSS 0
I_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VDDDM 1 AC=0.006944444444444444
V_X80Y20VDD_X80Y20VSS X80Y20VDDDM X80Y20VSS 0
I_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VDDDM 1 AC=0.006944444444444444
V_X80Y30VDD_X80Y30VSS X80Y30VDDDM X80Y30VSS 0
I_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VDDDM 1 AC=0.006944444444444444
V_X80Y40VDD_X80Y40VSS X80Y40VDDDM X80Y40VSS 0
I_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VDDDM 1 AC=0.006944444444444444
V_X80Y50VDD_X80Y50VSS X80Y50VDDDM X80Y50VSS 0
I_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VDDDM 1 AC=0.006944444444444444
V_X80Y60VDD_X80Y60VSS X80Y60VDDDM X80Y60VSS 0
I_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VDDDM 1 AC=0.006944444444444444
V_X80Y70VDD_X80Y70VSS X80Y70VDDDM X80Y70VSS 0
I_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VDDDM 1 AC=0.006944444444444444
V_X80Y80VDD_X80Y80VSS X80Y80VDDDM X80Y80VSS 0
I_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VDDDM 1 AC=0.006944444444444444
V_X80Y90VDD_X80Y90VSS X80Y90VDDDM X80Y90VSS 0
I_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VDDDM 1 AC=0.006944444444444444
V_X80Y100VDD_X80Y100VSS X80Y100VDDDM X80Y100VSS 0
I_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VDDDM 1 AC=0.006944444444444444
V_X80Y110VDD_X80Y110VSS X80Y110VDDDM X80Y110VSS 0
I_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VDDDM 1 AC=0.006944444444444444
V_X90Y120VDD_X90Y120VSS X90Y120VDDDM X90Y120VSS 0
I_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VDDDM 1 AC=0.006944444444444444
V_X90Y10VDD_X90Y10VSS X90Y10VDDDM X90Y10VSS 0
I_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VDDDM 1 AC=0.006944444444444444
V_X90Y20VDD_X90Y20VSS X90Y20VDDDM X90Y20VSS 0
I_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VDDDM 1 AC=0.006944444444444444
V_X90Y30VDD_X90Y30VSS X90Y30VDDDM X90Y30VSS 0
I_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VDDDM 1 AC=0.006944444444444444
V_X90Y40VDD_X90Y40VSS X90Y40VDDDM X90Y40VSS 0
I_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VDDDM 1 AC=0.006944444444444444
V_X90Y50VDD_X90Y50VSS X90Y50VDDDM X90Y50VSS 0
I_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VDDDM 1 AC=0.006944444444444444
V_X90Y60VDD_X90Y60VSS X90Y60VDDDM X90Y60VSS 0
I_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VDDDM 1 AC=0.006944444444444444
V_X90Y70VDD_X90Y70VSS X90Y70VDDDM X90Y70VSS 0
I_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VDDDM 1 AC=0.006944444444444444
V_X90Y80VDD_X90Y80VSS X90Y80VDDDM X90Y80VSS 0
I_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VDDDM 1 AC=0.006944444444444444
V_X90Y90VDD_X90Y90VSS X90Y90VDDDM X90Y90VSS 0
I_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VDDDM 1 AC=0.006944444444444444
V_X90Y100VDD_X90Y100VSS X90Y100VDDDM X90Y100VSS 0
I_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VDDDM 1 AC=0.006944444444444444
V_X90Y110VDD_X90Y110VSS X90Y110VDDDM X90Y110VSS 0
I_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VDDDM 1 AC=0.006944444444444444
V_X100Y120VDD_X100Y120VSS X100Y120VDDDM X100Y120VSS 0
I_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VDDDM 1 AC=0.006944444444444444
V_X100Y10VDD_X100Y10VSS X100Y10VDDDM X100Y10VSS 0
I_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VDDDM 1 AC=0.006944444444444444
V_X100Y20VDD_X100Y20VSS X100Y20VDDDM X100Y20VSS 0
I_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VDDDM 1 AC=0.006944444444444444
V_X100Y30VDD_X100Y30VSS X100Y30VDDDM X100Y30VSS 0
I_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VDDDM 1 AC=0.006944444444444444
V_X100Y40VDD_X100Y40VSS X100Y40VDDDM X100Y40VSS 0
I_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VDDDM 1 AC=0.006944444444444444
V_X100Y50VDD_X100Y50VSS X100Y50VDDDM X100Y50VSS 0
I_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VDDDM 1 AC=0.006944444444444444
V_X100Y60VDD_X100Y60VSS X100Y60VDDDM X100Y60VSS 0
I_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VDDDM 1 AC=0.006944444444444444
V_X100Y70VDD_X100Y70VSS X100Y70VDDDM X100Y70VSS 0
I_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VDDDM 1 AC=0.006944444444444444
V_X100Y80VDD_X100Y80VSS X100Y80VDDDM X100Y80VSS 0
I_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VDDDM 1 AC=0.006944444444444444
V_X100Y90VDD_X100Y90VSS X100Y90VDDDM X100Y90VSS 0
I_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VDDDM 1 AC=0.006944444444444444
V_X100Y100VDD_X100Y100VSS X100Y100VDDDM X100Y100VSS 0
I_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VDDDM 1 AC=0.006944444444444444
V_X100Y110VDD_X100Y110VSS X100Y110VDDDM X100Y110VSS 0
I_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VDDDM 1 AC=0.006944444444444444
V_X110Y120VDD_X110Y120VSS X110Y120VDDDM X110Y120VSS 0
I_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VDDDM 1 AC=0.006944444444444444
V_X110Y10VDD_X110Y10VSS X110Y10VDDDM X110Y10VSS 0
I_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VDDDM 1 AC=0.006944444444444444
V_X110Y20VDD_X110Y20VSS X110Y20VDDDM X110Y20VSS 0
I_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VDDDM 1 AC=0.006944444444444444
V_X110Y30VDD_X110Y30VSS X110Y30VDDDM X110Y30VSS 0
I_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VDDDM 1 AC=0.006944444444444444
V_X110Y40VDD_X110Y40VSS X110Y40VDDDM X110Y40VSS 0
I_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VDDDM 1 AC=0.006944444444444444
V_X110Y50VDD_X110Y50VSS X110Y50VDDDM X110Y50VSS 0
I_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VDDDM 1 AC=0.006944444444444444
V_X110Y60VDD_X110Y60VSS X110Y60VDDDM X110Y60VSS 0
I_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VDDDM 1 AC=0.006944444444444444
V_X110Y70VDD_X110Y70VSS X110Y70VDDDM X110Y70VSS 0
I_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VDDDM 1 AC=0.006944444444444444
V_X110Y80VDD_X110Y80VSS X110Y80VDDDM X110Y80VSS 0
I_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VDDDM 1 AC=0.006944444444444444
V_X110Y90VDD_X110Y90VSS X110Y90VDDDM X110Y90VSS 0
I_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VDDDM 1 AC=0.006944444444444444
V_X110Y100VDD_X110Y100VSS X110Y100VDDDM X110Y100VSS 0
I_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VDDDM 1 AC=0.006944444444444444
V_X110Y110VDD_X110Y110VSS X110Y110VDDDM X110Y110VSS 0
Rbump_X10Y10VDD X10Y10VDD X10Y10VDDM 20mOhm
Lbump_X10Y10VDD X10Y10VDDM VDD2 0.036nH
Rbump_X10Y10VSS X10Y10VSS X10Y10VSSM 20mOhm
Lbump_X10Y10VSS X10Y10VSSM VSS2 0.036nH
Rbump_X10Y20VDD X10Y20VDD X10Y20VDDM 20mOhm
Lbump_X10Y20VDD X10Y20VDDM VDD2 0.036nH
Rbump_X10Y20VSS X10Y20VSS X10Y20VSSM 20mOhm
Lbump_X10Y20VSS X10Y20VSSM VSS2 0.036nH
Rbump_X10Y30VDD X10Y30VDD X10Y30VDDM 20mOhm
Lbump_X10Y30VDD X10Y30VDDM VDD2 0.036nH
Rbump_X10Y30VSS X10Y30VSS X10Y30VSSM 20mOhm
Lbump_X10Y30VSS X10Y30VSSM VSS2 0.036nH
Rbump_X10Y40VDD X10Y40VDD X10Y40VDDM 20mOhm
Lbump_X10Y40VDD X10Y40VDDM VDD2 0.036nH
Rbump_X10Y40VSS X10Y40VSS X10Y40VSSM 20mOhm
Lbump_X10Y40VSS X10Y40VSSM VSS2 0.036nH
Rbump_X10Y50VDD X10Y50VDD X10Y50VDDM 20mOhm
Lbump_X10Y50VDD X10Y50VDDM VDD2 0.036nH
Rbump_X10Y50VSS X10Y50VSS X10Y50VSSM 20mOhm
Lbump_X10Y50VSS X10Y50VSSM VSS2 0.036nH
Rbump_X10Y60VDD X10Y60VDD X10Y60VDDM 20mOhm
Lbump_X10Y60VDD X10Y60VDDM VDD2 0.036nH
Rbump_X10Y60VSS X10Y60VSS X10Y60VSSM 20mOhm
Lbump_X10Y60VSS X10Y60VSSM VSS2 0.036nH
Rbump_X10Y70VDD X10Y70VDD X10Y70VDDM 20mOhm
Lbump_X10Y70VDD X10Y70VDDM VDD2 0.036nH
Rbump_X10Y70VSS X10Y70VSS X10Y70VSSM 20mOhm
Lbump_X10Y70VSS X10Y70VSSM VSS2 0.036nH
Rbump_X10Y80VDD X10Y80VDD X10Y80VDDM 20mOhm
Lbump_X10Y80VDD X10Y80VDDM VDD2 0.036nH
Rbump_X10Y80VSS X10Y80VSS X10Y80VSSM 20mOhm
Lbump_X10Y80VSS X10Y80VSSM VSS2 0.036nH
Rbump_X10Y90VDD X10Y90VDD X10Y90VDDM 20mOhm
Lbump_X10Y90VDD X10Y90VDDM VDD2 0.036nH
Rbump_X10Y90VSS X10Y90VSS X10Y90VSSM 20mOhm
Lbump_X10Y90VSS X10Y90VSSM VSS2 0.036nH
Rbump_X10Y100VDD X10Y100VDD X10Y100VDDM 20mOhm
Lbump_X10Y100VDD X10Y100VDDM VDD2 0.036nH
Rbump_X10Y100VSS X10Y100VSS X10Y100VSSM 20mOhm
Lbump_X10Y100VSS X10Y100VSSM VSS2 0.036nH
Rbump_X10Y110VDD X10Y110VDD X10Y110VDDM 20mOhm
Lbump_X10Y110VDD X10Y110VDDM VDD2 0.036nH
Rbump_X10Y110VSS X10Y110VSS X10Y110VSSM 20mOhm
Lbump_X10Y110VSS X10Y110VSSM VSS2 0.036nH
Rbump_X10Y120VDD X10Y120VDD X10Y120VDDM 20mOhm
Lbump_X10Y120VDD X10Y120VDDM VDD2 0.036nH
Rbump_X10Y120VSS X10Y120VSS X10Y120VSSM 20mOhm
Lbump_X10Y120VSS X10Y120VSSM VSS2 0.036nH
Rbump_X20Y10VDD X20Y10VDD X20Y10VDDM 20mOhm
Lbump_X20Y10VDD X20Y10VDDM VDD2 0.036nH
Rbump_X20Y10VSS X20Y10VSS X20Y10VSSM 20mOhm
Lbump_X20Y10VSS X20Y10VSSM VSS2 0.036nH
Rbump_X20Y20VDD X20Y20VDD X20Y20VDDM 20mOhm
Lbump_X20Y20VDD X20Y20VDDM VDD2 0.036nH
Rbump_X20Y20VSS X20Y20VSS X20Y20VSSM 20mOhm
Lbump_X20Y20VSS X20Y20VSSM VSS2 0.036nH
Rbump_X20Y30VDD X20Y30VDD X20Y30VDDM 20mOhm
Lbump_X20Y30VDD X20Y30VDDM VDD2 0.036nH
Rbump_X20Y30VSS X20Y30VSS X20Y30VSSM 20mOhm
Lbump_X20Y30VSS X20Y30VSSM VSS2 0.036nH
Rbump_X20Y40VDD X20Y40VDD X20Y40VDDM 20mOhm
Lbump_X20Y40VDD X20Y40VDDM VDD2 0.036nH
Rbump_X20Y40VSS X20Y40VSS X20Y40VSSM 20mOhm
Lbump_X20Y40VSS X20Y40VSSM VSS2 0.036nH
Rbump_X20Y50VDD X20Y50VDD X20Y50VDDM 20mOhm
Lbump_X20Y50VDD X20Y50VDDM VDD2 0.036nH
Rbump_X20Y50VSS X20Y50VSS X20Y50VSSM 20mOhm
Lbump_X20Y50VSS X20Y50VSSM VSS2 0.036nH
Rbump_X20Y60VDD X20Y60VDD X20Y60VDDM 20mOhm
Lbump_X20Y60VDD X20Y60VDDM VDD2 0.036nH
Rbump_X20Y60VSS X20Y60VSS X20Y60VSSM 20mOhm
Lbump_X20Y60VSS X20Y60VSSM VSS2 0.036nH
Rbump_X20Y70VDD X20Y70VDD X20Y70VDDM 20mOhm
Lbump_X20Y70VDD X20Y70VDDM VDD2 0.036nH
Rbump_X20Y70VSS X20Y70VSS X20Y70VSSM 20mOhm
Lbump_X20Y70VSS X20Y70VSSM VSS2 0.036nH
Rbump_X20Y80VDD X20Y80VDD X20Y80VDDM 20mOhm
Lbump_X20Y80VDD X20Y80VDDM VDD2 0.036nH
Rbump_X20Y80VSS X20Y80VSS X20Y80VSSM 20mOhm
Lbump_X20Y80VSS X20Y80VSSM VSS2 0.036nH
Rbump_X20Y90VDD X20Y90VDD X20Y90VDDM 20mOhm
Lbump_X20Y90VDD X20Y90VDDM VDD2 0.036nH
Rbump_X20Y90VSS X20Y90VSS X20Y90VSSM 20mOhm
Lbump_X20Y90VSS X20Y90VSSM VSS2 0.036nH
Rbump_X20Y100VDD X20Y100VDD X20Y100VDDM 20mOhm
Lbump_X20Y100VDD X20Y100VDDM VDD2 0.036nH
Rbump_X20Y100VSS X20Y100VSS X20Y100VSSM 20mOhm
Lbump_X20Y100VSS X20Y100VSSM VSS2 0.036nH
Rbump_X20Y110VDD X20Y110VDD X20Y110VDDM 20mOhm
Lbump_X20Y110VDD X20Y110VDDM VDD2 0.036nH
Rbump_X20Y110VSS X20Y110VSS X20Y110VSSM 20mOhm
Lbump_X20Y110VSS X20Y110VSSM VSS2 0.036nH
Rbump_X20Y120VDD X20Y120VDD X20Y120VDDM 20mOhm
Lbump_X20Y120VDD X20Y120VDDM VDD2 0.036nH
Rbump_X20Y120VSS X20Y120VSS X20Y120VSSM 20mOhm
Lbump_X20Y120VSS X20Y120VSSM VSS2 0.036nH
Rbump_X30Y10VDD X30Y10VDD X30Y10VDDM 20mOhm
Lbump_X30Y10VDD X30Y10VDDM VDD2 0.036nH
Rbump_X30Y10VSS X30Y10VSS X30Y10VSSM 20mOhm
Lbump_X30Y10VSS X30Y10VSSM VSS2 0.036nH
Rbump_X30Y20VDD X30Y20VDD X30Y20VDDM 20mOhm
Lbump_X30Y20VDD X30Y20VDDM VDD2 0.036nH
Rbump_X30Y20VSS X30Y20VSS X30Y20VSSM 20mOhm
Lbump_X30Y20VSS X30Y20VSSM VSS2 0.036nH
Rbump_X30Y30VDD X30Y30VDD X30Y30VDDM 20mOhm
Lbump_X30Y30VDD X30Y30VDDM VDD2 0.036nH
Rbump_X30Y30VSS X30Y30VSS X30Y30VSSM 20mOhm
Lbump_X30Y30VSS X30Y30VSSM VSS2 0.036nH
Rbump_X30Y40VDD X30Y40VDD X30Y40VDDM 20mOhm
Lbump_X30Y40VDD X30Y40VDDM VDD2 0.036nH
Rbump_X30Y40VSS X30Y40VSS X30Y40VSSM 20mOhm
Lbump_X30Y40VSS X30Y40VSSM VSS2 0.036nH
Rbump_X30Y50VDD X30Y50VDD X30Y50VDDM 20mOhm
Lbump_X30Y50VDD X30Y50VDDM VDD2 0.036nH
Rbump_X30Y50VSS X30Y50VSS X30Y50VSSM 20mOhm
Lbump_X30Y50VSS X30Y50VSSM VSS2 0.036nH
Rbump_X30Y60VDD X30Y60VDD X30Y60VDDM 20mOhm
Lbump_X30Y60VDD X30Y60VDDM VDD2 0.036nH
Rbump_X30Y60VSS X30Y60VSS X30Y60VSSM 20mOhm
Lbump_X30Y60VSS X30Y60VSSM VSS2 0.036nH
Rbump_X30Y70VDD X30Y70VDD X30Y70VDDM 20mOhm
Lbump_X30Y70VDD X30Y70VDDM VDD2 0.036nH
Rbump_X30Y70VSS X30Y70VSS X30Y70VSSM 20mOhm
Lbump_X30Y70VSS X30Y70VSSM VSS2 0.036nH
Rbump_X30Y80VDD X30Y80VDD X30Y80VDDM 20mOhm
Lbump_X30Y80VDD X30Y80VDDM VDD2 0.036nH
Rbump_X30Y80VSS X30Y80VSS X30Y80VSSM 20mOhm
Lbump_X30Y80VSS X30Y80VSSM VSS2 0.036nH
Rbump_X30Y90VDD X30Y90VDD X30Y90VDDM 20mOhm
Lbump_X30Y90VDD X30Y90VDDM VDD2 0.036nH
Rbump_X30Y90VSS X30Y90VSS X30Y90VSSM 20mOhm
Lbump_X30Y90VSS X30Y90VSSM VSS2 0.036nH
Rbump_X30Y100VDD X30Y100VDD X30Y100VDDM 20mOhm
Lbump_X30Y100VDD X30Y100VDDM VDD2 0.036nH
Rbump_X30Y100VSS X30Y100VSS X30Y100VSSM 20mOhm
Lbump_X30Y100VSS X30Y100VSSM VSS2 0.036nH
Rbump_X30Y110VDD X30Y110VDD X30Y110VDDM 20mOhm
Lbump_X30Y110VDD X30Y110VDDM VDD2 0.036nH
Rbump_X30Y110VSS X30Y110VSS X30Y110VSSM 20mOhm
Lbump_X30Y110VSS X30Y110VSSM VSS2 0.036nH
Rbump_X30Y120VDD X30Y120VDD X30Y120VDDM 20mOhm
Lbump_X30Y120VDD X30Y120VDDM VDD2 0.036nH
Rbump_X30Y120VSS X30Y120VSS X30Y120VSSM 20mOhm
Lbump_X30Y120VSS X30Y120VSSM VSS2 0.036nH
Rbump_X40Y10VDD X40Y10VDD X40Y10VDDM 20mOhm
Lbump_X40Y10VDD X40Y10VDDM VDD2 0.036nH
Rbump_X40Y10VSS X40Y10VSS X40Y10VSSM 20mOhm
Lbump_X40Y10VSS X40Y10VSSM VSS2 0.036nH
Rbump_X40Y20VDD X40Y20VDD X40Y20VDDM 20mOhm
Lbump_X40Y20VDD X40Y20VDDM VDD2 0.036nH
Rbump_X40Y20VSS X40Y20VSS X40Y20VSSM 20mOhm
Lbump_X40Y20VSS X40Y20VSSM VSS2 0.036nH
Rbump_X40Y30VDD X40Y30VDD X40Y30VDDM 20mOhm
Lbump_X40Y30VDD X40Y30VDDM VDD2 0.036nH
Rbump_X40Y30VSS X40Y30VSS X40Y30VSSM 20mOhm
Lbump_X40Y30VSS X40Y30VSSM VSS2 0.036nH
Rbump_X40Y40VDD X40Y40VDD X40Y40VDDM 20mOhm
Lbump_X40Y40VDD X40Y40VDDM VDD2 0.036nH
Rbump_X40Y40VSS X40Y40VSS X40Y40VSSM 20mOhm
Lbump_X40Y40VSS X40Y40VSSM VSS2 0.036nH
Rbump_X40Y50VDD X40Y50VDD X40Y50VDDM 20mOhm
Lbump_X40Y50VDD X40Y50VDDM VDD2 0.036nH
Rbump_X40Y50VSS X40Y50VSS X40Y50VSSM 20mOhm
Lbump_X40Y50VSS X40Y50VSSM VSS2 0.036nH
Rbump_X40Y60VDD X40Y60VDD X40Y60VDDM 20mOhm
Lbump_X40Y60VDD X40Y60VDDM VDD2 0.036nH
Rbump_X40Y60VSS X40Y60VSS X40Y60VSSM 20mOhm
Lbump_X40Y60VSS X40Y60VSSM VSS2 0.036nH
Rbump_X40Y70VDD X40Y70VDD X40Y70VDDM 20mOhm
Lbump_X40Y70VDD X40Y70VDDM VDD2 0.036nH
Rbump_X40Y70VSS X40Y70VSS X40Y70VSSM 20mOhm
Lbump_X40Y70VSS X40Y70VSSM VSS2 0.036nH
Rbump_X40Y80VDD X40Y80VDD X40Y80VDDM 20mOhm
Lbump_X40Y80VDD X40Y80VDDM VDD2 0.036nH
Rbump_X40Y80VSS X40Y80VSS X40Y80VSSM 20mOhm
Lbump_X40Y80VSS X40Y80VSSM VSS2 0.036nH
Rbump_X40Y90VDD X40Y90VDD X40Y90VDDM 20mOhm
Lbump_X40Y90VDD X40Y90VDDM VDD2 0.036nH
Rbump_X40Y90VSS X40Y90VSS X40Y90VSSM 20mOhm
Lbump_X40Y90VSS X40Y90VSSM VSS2 0.036nH
Rbump_X40Y100VDD X40Y100VDD X40Y100VDDM 20mOhm
Lbump_X40Y100VDD X40Y100VDDM VDD2 0.036nH
Rbump_X40Y100VSS X40Y100VSS X40Y100VSSM 20mOhm
Lbump_X40Y100VSS X40Y100VSSM VSS2 0.036nH
Rbump_X40Y110VDD X40Y110VDD X40Y110VDDM 20mOhm
Lbump_X40Y110VDD X40Y110VDDM VDD2 0.036nH
Rbump_X40Y110VSS X40Y110VSS X40Y110VSSM 20mOhm
Lbump_X40Y110VSS X40Y110VSSM VSS2 0.036nH
Rbump_X40Y120VDD X40Y120VDD X40Y120VDDM 20mOhm
Lbump_X40Y120VDD X40Y120VDDM VDD2 0.036nH
Rbump_X40Y120VSS X40Y120VSS X40Y120VSSM 20mOhm
Lbump_X40Y120VSS X40Y120VSSM VSS2 0.036nH
Rbump_X50Y10VDD X50Y10VDD X50Y10VDDM 20mOhm
Lbump_X50Y10VDD X50Y10VDDM VDD2 0.036nH
Rbump_X50Y10VSS X50Y10VSS X50Y10VSSM 20mOhm
Lbump_X50Y10VSS X50Y10VSSM VSS2 0.036nH
Rbump_X50Y20VDD X50Y20VDD X50Y20VDDM 20mOhm
Lbump_X50Y20VDD X50Y20VDDM VDD2 0.036nH
Rbump_X50Y20VSS X50Y20VSS X50Y20VSSM 20mOhm
Lbump_X50Y20VSS X50Y20VSSM VSS2 0.036nH
Rbump_X50Y30VDD X50Y30VDD X50Y30VDDM 20mOhm
Lbump_X50Y30VDD X50Y30VDDM VDD2 0.036nH
Rbump_X50Y30VSS X50Y30VSS X50Y30VSSM 20mOhm
Lbump_X50Y30VSS X50Y30VSSM VSS2 0.036nH
Rbump_X50Y40VDD X50Y40VDD X50Y40VDDM 20mOhm
Lbump_X50Y40VDD X50Y40VDDM VDD2 0.036nH
Rbump_X50Y40VSS X50Y40VSS X50Y40VSSM 20mOhm
Lbump_X50Y40VSS X50Y40VSSM VSS2 0.036nH
Rbump_X50Y50VDD X50Y50VDD X50Y50VDDM 20mOhm
Lbump_X50Y50VDD X50Y50VDDM VDD2 0.036nH
Rbump_X50Y50VSS X50Y50VSS X50Y50VSSM 20mOhm
Lbump_X50Y50VSS X50Y50VSSM VSS2 0.036nH
Rbump_X50Y60VDD X50Y60VDD X50Y60VDDM 20mOhm
Lbump_X50Y60VDD X50Y60VDDM VDD2 0.036nH
Rbump_X50Y60VSS X50Y60VSS X50Y60VSSM 20mOhm
Lbump_X50Y60VSS X50Y60VSSM VSS2 0.036nH
Rbump_X50Y70VDD X50Y70VDD X50Y70VDDM 20mOhm
Lbump_X50Y70VDD X50Y70VDDM VDD2 0.036nH
Rbump_X50Y70VSS X50Y70VSS X50Y70VSSM 20mOhm
Lbump_X50Y70VSS X50Y70VSSM VSS2 0.036nH
Rbump_X50Y80VDD X50Y80VDD X50Y80VDDM 20mOhm
Lbump_X50Y80VDD X50Y80VDDM VDD2 0.036nH
Rbump_X50Y80VSS X50Y80VSS X50Y80VSSM 20mOhm
Lbump_X50Y80VSS X50Y80VSSM VSS2 0.036nH
Rbump_X50Y90VDD X50Y90VDD X50Y90VDDM 20mOhm
Lbump_X50Y90VDD X50Y90VDDM VDD2 0.036nH
Rbump_X50Y90VSS X50Y90VSS X50Y90VSSM 20mOhm
Lbump_X50Y90VSS X50Y90VSSM VSS2 0.036nH
Rbump_X50Y100VDD X50Y100VDD X50Y100VDDM 20mOhm
Lbump_X50Y100VDD X50Y100VDDM VDD2 0.036nH
Rbump_X50Y100VSS X50Y100VSS X50Y100VSSM 20mOhm
Lbump_X50Y100VSS X50Y100VSSM VSS2 0.036nH
Rbump_X50Y110VDD X50Y110VDD X50Y110VDDM 20mOhm
Lbump_X50Y110VDD X50Y110VDDM VDD2 0.036nH
Rbump_X50Y110VSS X50Y110VSS X50Y110VSSM 20mOhm
Lbump_X50Y110VSS X50Y110VSSM VSS2 0.036nH
Rbump_X50Y120VDD X50Y120VDD X50Y120VDDM 20mOhm
Lbump_X50Y120VDD X50Y120VDDM VDD2 0.036nH
Rbump_X50Y120VSS X50Y120VSS X50Y120VSSM 20mOhm
Lbump_X50Y120VSS X50Y120VSSM VSS2 0.036nH
Rbump_X60Y10VDD X60Y10VDD X60Y10VDDM 20mOhm
Lbump_X60Y10VDD X60Y10VDDM VDD2 0.036nH
Rbump_X60Y10VSS X60Y10VSS X60Y10VSSM 20mOhm
Lbump_X60Y10VSS X60Y10VSSM VSS2 0.036nH
Rbump_X60Y20VDD X60Y20VDD X60Y20VDDM 20mOhm
Lbump_X60Y20VDD X60Y20VDDM VDD2 0.036nH
Rbump_X60Y20VSS X60Y20VSS X60Y20VSSM 20mOhm
Lbump_X60Y20VSS X60Y20VSSM VSS2 0.036nH
Rbump_X60Y30VDD X60Y30VDD X60Y30VDDM 20mOhm
Lbump_X60Y30VDD X60Y30VDDM VDD2 0.036nH
Rbump_X60Y30VSS X60Y30VSS X60Y30VSSM 20mOhm
Lbump_X60Y30VSS X60Y30VSSM VSS2 0.036nH
Rbump_X60Y40VDD X60Y40VDD X60Y40VDDM 20mOhm
Lbump_X60Y40VDD X60Y40VDDM VDD2 0.036nH
Rbump_X60Y40VSS X60Y40VSS X60Y40VSSM 20mOhm
Lbump_X60Y40VSS X60Y40VSSM VSS2 0.036nH
Rbump_X60Y50VDD X60Y50VDD X60Y50VDDM 20mOhm
Lbump_X60Y50VDD X60Y50VDDM VDD2 0.036nH
Rbump_X60Y50VSS X60Y50VSS X60Y50VSSM 20mOhm
Lbump_X60Y50VSS X60Y50VSSM VSS2 0.036nH
Rbump_X60Y60VDD X60Y60VDD X60Y60VDDM 20mOhm
Lbump_X60Y60VDD X60Y60VDDM VDD2 0.036nH
Rbump_X60Y60VSS X60Y60VSS X60Y60VSSM 20mOhm
Lbump_X60Y60VSS X60Y60VSSM VSS2 0.036nH
Rbump_X60Y70VDD X60Y70VDD X60Y70VDDM 20mOhm
Lbump_X60Y70VDD X60Y70VDDM VDD2 0.036nH
Rbump_X60Y70VSS X60Y70VSS X60Y70VSSM 20mOhm
Lbump_X60Y70VSS X60Y70VSSM VSS2 0.036nH
Rbump_X60Y80VDD X60Y80VDD X60Y80VDDM 20mOhm
Lbump_X60Y80VDD X60Y80VDDM VDD2 0.036nH
Rbump_X60Y80VSS X60Y80VSS X60Y80VSSM 20mOhm
Lbump_X60Y80VSS X60Y80VSSM VSS2 0.036nH
Rbump_X60Y90VDD X60Y90VDD X60Y90VDDM 20mOhm
Lbump_X60Y90VDD X60Y90VDDM VDD2 0.036nH
Rbump_X60Y90VSS X60Y90VSS X60Y90VSSM 20mOhm
Lbump_X60Y90VSS X60Y90VSSM VSS2 0.036nH
Rbump_X60Y100VDD X60Y100VDD X60Y100VDDM 20mOhm
Lbump_X60Y100VDD X60Y100VDDM VDD2 0.036nH
Rbump_X60Y100VSS X60Y100VSS X60Y100VSSM 20mOhm
Lbump_X60Y100VSS X60Y100VSSM VSS2 0.036nH
Rbump_X60Y110VDD X60Y110VDD X60Y110VDDM 20mOhm
Lbump_X60Y110VDD X60Y110VDDM VDD2 0.036nH
Rbump_X60Y110VSS X60Y110VSS X60Y110VSSM 20mOhm
Lbump_X60Y110VSS X60Y110VSSM VSS2 0.036nH
Rbump_X60Y120VDD X60Y120VDD X60Y120VDDM 20mOhm
Lbump_X60Y120VDD X60Y120VDDM VDD2 0.036nH
Rbump_X60Y120VSS X60Y120VSS X60Y120VSSM 20mOhm
Lbump_X60Y120VSS X60Y120VSSM VSS2 0.036nH
Rbump_X70Y10VDD X70Y10VDD X70Y10VDDM 20mOhm
Lbump_X70Y10VDD X70Y10VDDM VDD2 0.036nH
Rbump_X70Y10VSS X70Y10VSS X70Y10VSSM 20mOhm
Lbump_X70Y10VSS X70Y10VSSM VSS2 0.036nH
Rbump_X70Y20VDD X70Y20VDD X70Y20VDDM 20mOhm
Lbump_X70Y20VDD X70Y20VDDM VDD2 0.036nH
Rbump_X70Y20VSS X70Y20VSS X70Y20VSSM 20mOhm
Lbump_X70Y20VSS X70Y20VSSM VSS2 0.036nH
Rbump_X70Y30VDD X70Y30VDD X70Y30VDDM 20mOhm
Lbump_X70Y30VDD X70Y30VDDM VDD2 0.036nH
Rbump_X70Y30VSS X70Y30VSS X70Y30VSSM 20mOhm
Lbump_X70Y30VSS X70Y30VSSM VSS2 0.036nH
Rbump_X70Y40VDD X70Y40VDD X70Y40VDDM 20mOhm
Lbump_X70Y40VDD X70Y40VDDM VDD2 0.036nH
Rbump_X70Y40VSS X70Y40VSS X70Y40VSSM 20mOhm
Lbump_X70Y40VSS X70Y40VSSM VSS2 0.036nH
Rbump_X70Y50VDD X70Y50VDD X70Y50VDDM 20mOhm
Lbump_X70Y50VDD X70Y50VDDM VDD2 0.036nH
Rbump_X70Y50VSS X70Y50VSS X70Y50VSSM 20mOhm
Lbump_X70Y50VSS X70Y50VSSM VSS2 0.036nH
Rbump_X70Y60VDD X70Y60VDD X70Y60VDDM 20mOhm
Lbump_X70Y60VDD X70Y60VDDM VDD2 0.036nH
Rbump_X70Y60VSS X70Y60VSS X70Y60VSSM 20mOhm
Lbump_X70Y60VSS X70Y60VSSM VSS2 0.036nH
Rbump_X70Y70VDD X70Y70VDD X70Y70VDDM 20mOhm
Lbump_X70Y70VDD X70Y70VDDM VDD2 0.036nH
Rbump_X70Y70VSS X70Y70VSS X70Y70VSSM 20mOhm
Lbump_X70Y70VSS X70Y70VSSM VSS2 0.036nH
Rbump_X70Y80VDD X70Y80VDD X70Y80VDDM 20mOhm
Lbump_X70Y80VDD X70Y80VDDM VDD2 0.036nH
Rbump_X70Y80VSS X70Y80VSS X70Y80VSSM 20mOhm
Lbump_X70Y80VSS X70Y80VSSM VSS2 0.036nH
Rbump_X70Y90VDD X70Y90VDD X70Y90VDDM 20mOhm
Lbump_X70Y90VDD X70Y90VDDM VDD2 0.036nH
Rbump_X70Y90VSS X70Y90VSS X70Y90VSSM 20mOhm
Lbump_X70Y90VSS X70Y90VSSM VSS2 0.036nH
Rbump_X70Y100VDD X70Y100VDD X70Y100VDDM 20mOhm
Lbump_X70Y100VDD X70Y100VDDM VDD2 0.036nH
Rbump_X70Y100VSS X70Y100VSS X70Y100VSSM 20mOhm
Lbump_X70Y100VSS X70Y100VSSM VSS2 0.036nH
Rbump_X70Y110VDD X70Y110VDD X70Y110VDDM 20mOhm
Lbump_X70Y110VDD X70Y110VDDM VDD2 0.036nH
Rbump_X70Y110VSS X70Y110VSS X70Y110VSSM 20mOhm
Lbump_X70Y110VSS X70Y110VSSM VSS2 0.036nH
Rbump_X70Y120VDD X70Y120VDD X70Y120VDDM 20mOhm
Lbump_X70Y120VDD X70Y120VDDM VDD2 0.036nH
Rbump_X70Y120VSS X70Y120VSS X70Y120VSSM 20mOhm
Lbump_X70Y120VSS X70Y120VSSM VSS2 0.036nH
Rbump_X80Y10VDD X80Y10VDD X80Y10VDDM 20mOhm
Lbump_X80Y10VDD X80Y10VDDM VDD2 0.036nH
Rbump_X80Y10VSS X80Y10VSS X80Y10VSSM 20mOhm
Lbump_X80Y10VSS X80Y10VSSM VSS2 0.036nH
Rbump_X80Y20VDD X80Y20VDD X80Y20VDDM 20mOhm
Lbump_X80Y20VDD X80Y20VDDM VDD2 0.036nH
Rbump_X80Y20VSS X80Y20VSS X80Y20VSSM 20mOhm
Lbump_X80Y20VSS X80Y20VSSM VSS2 0.036nH
Rbump_X80Y30VDD X80Y30VDD X80Y30VDDM 20mOhm
Lbump_X80Y30VDD X80Y30VDDM VDD2 0.036nH
Rbump_X80Y30VSS X80Y30VSS X80Y30VSSM 20mOhm
Lbump_X80Y30VSS X80Y30VSSM VSS2 0.036nH
Rbump_X80Y40VDD X80Y40VDD X80Y40VDDM 20mOhm
Lbump_X80Y40VDD X80Y40VDDM VDD2 0.036nH
Rbump_X80Y40VSS X80Y40VSS X80Y40VSSM 20mOhm
Lbump_X80Y40VSS X80Y40VSSM VSS2 0.036nH
Rbump_X80Y50VDD X80Y50VDD X80Y50VDDM 20mOhm
Lbump_X80Y50VDD X80Y50VDDM VDD2 0.036nH
Rbump_X80Y50VSS X80Y50VSS X80Y50VSSM 20mOhm
Lbump_X80Y50VSS X80Y50VSSM VSS2 0.036nH
Rbump_X80Y60VDD X80Y60VDD X80Y60VDDM 20mOhm
Lbump_X80Y60VDD X80Y60VDDM VDD2 0.036nH
Rbump_X80Y60VSS X80Y60VSS X80Y60VSSM 20mOhm
Lbump_X80Y60VSS X80Y60VSSM VSS2 0.036nH
Rbump_X80Y70VDD X80Y70VDD X80Y70VDDM 20mOhm
Lbump_X80Y70VDD X80Y70VDDM VDD2 0.036nH
Rbump_X80Y70VSS X80Y70VSS X80Y70VSSM 20mOhm
Lbump_X80Y70VSS X80Y70VSSM VSS2 0.036nH
Rbump_X80Y80VDD X80Y80VDD X80Y80VDDM 20mOhm
Lbump_X80Y80VDD X80Y80VDDM VDD2 0.036nH
Rbump_X80Y80VSS X80Y80VSS X80Y80VSSM 20mOhm
Lbump_X80Y80VSS X80Y80VSSM VSS2 0.036nH
Rbump_X80Y90VDD X80Y90VDD X80Y90VDDM 20mOhm
Lbump_X80Y90VDD X80Y90VDDM VDD2 0.036nH
Rbump_X80Y90VSS X80Y90VSS X80Y90VSSM 20mOhm
Lbump_X80Y90VSS X80Y90VSSM VSS2 0.036nH
Rbump_X80Y100VDD X80Y100VDD X80Y100VDDM 20mOhm
Lbump_X80Y100VDD X80Y100VDDM VDD2 0.036nH
Rbump_X80Y100VSS X80Y100VSS X80Y100VSSM 20mOhm
Lbump_X80Y100VSS X80Y100VSSM VSS2 0.036nH
Rbump_X80Y110VDD X80Y110VDD X80Y110VDDM 20mOhm
Lbump_X80Y110VDD X80Y110VDDM VDD2 0.036nH
Rbump_X80Y110VSS X80Y110VSS X80Y110VSSM 20mOhm
Lbump_X80Y110VSS X80Y110VSSM VSS2 0.036nH
Rbump_X80Y120VDD X80Y120VDD X80Y120VDDM 20mOhm
Lbump_X80Y120VDD X80Y120VDDM VDD2 0.036nH
Rbump_X80Y120VSS X80Y120VSS X80Y120VSSM 20mOhm
Lbump_X80Y120VSS X80Y120VSSM VSS2 0.036nH
Rbump_X90Y10VDD X90Y10VDD X90Y10VDDM 20mOhm
Lbump_X90Y10VDD X90Y10VDDM VDD2 0.036nH
Rbump_X90Y10VSS X90Y10VSS X90Y10VSSM 20mOhm
Lbump_X90Y10VSS X90Y10VSSM VSS2 0.036nH
Rbump_X90Y20VDD X90Y20VDD X90Y20VDDM 20mOhm
Lbump_X90Y20VDD X90Y20VDDM VDD2 0.036nH
Rbump_X90Y20VSS X90Y20VSS X90Y20VSSM 20mOhm
Lbump_X90Y20VSS X90Y20VSSM VSS2 0.036nH
Rbump_X90Y30VDD X90Y30VDD X90Y30VDDM 20mOhm
Lbump_X90Y30VDD X90Y30VDDM VDD2 0.036nH
Rbump_X90Y30VSS X90Y30VSS X90Y30VSSM 20mOhm
Lbump_X90Y30VSS X90Y30VSSM VSS2 0.036nH
Rbump_X90Y40VDD X90Y40VDD X90Y40VDDM 20mOhm
Lbump_X90Y40VDD X90Y40VDDM VDD2 0.036nH
Rbump_X90Y40VSS X90Y40VSS X90Y40VSSM 20mOhm
Lbump_X90Y40VSS X90Y40VSSM VSS2 0.036nH
Rbump_X90Y50VDD X90Y50VDD X90Y50VDDM 20mOhm
Lbump_X90Y50VDD X90Y50VDDM VDD2 0.036nH
Rbump_X90Y50VSS X90Y50VSS X90Y50VSSM 20mOhm
Lbump_X90Y50VSS X90Y50VSSM VSS2 0.036nH
Rbump_X90Y60VDD X90Y60VDD X90Y60VDDM 20mOhm
Lbump_X90Y60VDD X90Y60VDDM VDD2 0.036nH
Rbump_X90Y60VSS X90Y60VSS X90Y60VSSM 20mOhm
Lbump_X90Y60VSS X90Y60VSSM VSS2 0.036nH
Rbump_X90Y70VDD X90Y70VDD X90Y70VDDM 20mOhm
Lbump_X90Y70VDD X90Y70VDDM VDD2 0.036nH
Rbump_X90Y70VSS X90Y70VSS X90Y70VSSM 20mOhm
Lbump_X90Y70VSS X90Y70VSSM VSS2 0.036nH
Rbump_X90Y80VDD X90Y80VDD X90Y80VDDM 20mOhm
Lbump_X90Y80VDD X90Y80VDDM VDD2 0.036nH
Rbump_X90Y80VSS X90Y80VSS X90Y80VSSM 20mOhm
Lbump_X90Y80VSS X90Y80VSSM VSS2 0.036nH
Rbump_X90Y90VDD X90Y90VDD X90Y90VDDM 20mOhm
Lbump_X90Y90VDD X90Y90VDDM VDD2 0.036nH
Rbump_X90Y90VSS X90Y90VSS X90Y90VSSM 20mOhm
Lbump_X90Y90VSS X90Y90VSSM VSS2 0.036nH
Rbump_X90Y100VDD X90Y100VDD X90Y100VDDM 20mOhm
Lbump_X90Y100VDD X90Y100VDDM VDD2 0.036nH
Rbump_X90Y100VSS X90Y100VSS X90Y100VSSM 20mOhm
Lbump_X90Y100VSS X90Y100VSSM VSS2 0.036nH
Rbump_X90Y110VDD X90Y110VDD X90Y110VDDM 20mOhm
Lbump_X90Y110VDD X90Y110VDDM VDD2 0.036nH
Rbump_X90Y110VSS X90Y110VSS X90Y110VSSM 20mOhm
Lbump_X90Y110VSS X90Y110VSSM VSS2 0.036nH
Rbump_X90Y120VDD X90Y120VDD X90Y120VDDM 20mOhm
Lbump_X90Y120VDD X90Y120VDDM VDD2 0.036nH
Rbump_X90Y120VSS X90Y120VSS X90Y120VSSM 20mOhm
Lbump_X90Y120VSS X90Y120VSSM VSS2 0.036nH
Rbump_X100Y10VDD X100Y10VDD X100Y10VDDM 20mOhm
Lbump_X100Y10VDD X100Y10VDDM VDD2 0.036nH
Rbump_X100Y10VSS X100Y10VSS X100Y10VSSM 20mOhm
Lbump_X100Y10VSS X100Y10VSSM VSS2 0.036nH
Rbump_X100Y20VDD X100Y20VDD X100Y20VDDM 20mOhm
Lbump_X100Y20VDD X100Y20VDDM VDD2 0.036nH
Rbump_X100Y20VSS X100Y20VSS X100Y20VSSM 20mOhm
Lbump_X100Y20VSS X100Y20VSSM VSS2 0.036nH
Rbump_X100Y30VDD X100Y30VDD X100Y30VDDM 20mOhm
Lbump_X100Y30VDD X100Y30VDDM VDD2 0.036nH
Rbump_X100Y30VSS X100Y30VSS X100Y30VSSM 20mOhm
Lbump_X100Y30VSS X100Y30VSSM VSS2 0.036nH
Rbump_X100Y40VDD X100Y40VDD X100Y40VDDM 20mOhm
Lbump_X100Y40VDD X100Y40VDDM VDD2 0.036nH
Rbump_X100Y40VSS X100Y40VSS X100Y40VSSM 20mOhm
Lbump_X100Y40VSS X100Y40VSSM VSS2 0.036nH
Rbump_X100Y50VDD X100Y50VDD X100Y50VDDM 20mOhm
Lbump_X100Y50VDD X100Y50VDDM VDD2 0.036nH
Rbump_X100Y50VSS X100Y50VSS X100Y50VSSM 20mOhm
Lbump_X100Y50VSS X100Y50VSSM VSS2 0.036nH
Rbump_X100Y60VDD X100Y60VDD X100Y60VDDM 20mOhm
Lbump_X100Y60VDD X100Y60VDDM VDD2 0.036nH
Rbump_X100Y60VSS X100Y60VSS X100Y60VSSM 20mOhm
Lbump_X100Y60VSS X100Y60VSSM VSS2 0.036nH
Rbump_X100Y70VDD X100Y70VDD X100Y70VDDM 20mOhm
Lbump_X100Y70VDD X100Y70VDDM VDD2 0.036nH
Rbump_X100Y70VSS X100Y70VSS X100Y70VSSM 20mOhm
Lbump_X100Y70VSS X100Y70VSSM VSS2 0.036nH
Rbump_X100Y80VDD X100Y80VDD X100Y80VDDM 20mOhm
Lbump_X100Y80VDD X100Y80VDDM VDD2 0.036nH
Rbump_X100Y80VSS X100Y80VSS X100Y80VSSM 20mOhm
Lbump_X100Y80VSS X100Y80VSSM VSS2 0.036nH
Rbump_X100Y90VDD X100Y90VDD X100Y90VDDM 20mOhm
Lbump_X100Y90VDD X100Y90VDDM VDD2 0.036nH
Rbump_X100Y90VSS X100Y90VSS X100Y90VSSM 20mOhm
Lbump_X100Y90VSS X100Y90VSSM VSS2 0.036nH
Rbump_X100Y100VDD X100Y100VDD X100Y100VDDM 20mOhm
Lbump_X100Y100VDD X100Y100VDDM VDD2 0.036nH
Rbump_X100Y100VSS X100Y100VSS X100Y100VSSM 20mOhm
Lbump_X100Y100VSS X100Y100VSSM VSS2 0.036nH
Rbump_X100Y110VDD X100Y110VDD X100Y110VDDM 20mOhm
Lbump_X100Y110VDD X100Y110VDDM VDD2 0.036nH
Rbump_X100Y110VSS X100Y110VSS X100Y110VSSM 20mOhm
Lbump_X100Y110VSS X100Y110VSSM VSS2 0.036nH
Rbump_X100Y120VDD X100Y120VDD X100Y120VDDM 20mOhm
Lbump_X100Y120VDD X100Y120VDDM VDD2 0.036nH
Rbump_X100Y120VSS X100Y120VSS X100Y120VSSM 20mOhm
Lbump_X100Y120VSS X100Y120VSSM VSS2 0.036nH
Rbump_X110Y10VDD X110Y10VDD X110Y10VDDM 20mOhm
Lbump_X110Y10VDD X110Y10VDDM VDD2 0.036nH
Rbump_X110Y10VSS X110Y10VSS X110Y10VSSM 20mOhm
Lbump_X110Y10VSS X110Y10VSSM VSS2 0.036nH
Rbump_X110Y20VDD X110Y20VDD X110Y20VDDM 20mOhm
Lbump_X110Y20VDD X110Y20VDDM VDD2 0.036nH
Rbump_X110Y20VSS X110Y20VSS X110Y20VSSM 20mOhm
Lbump_X110Y20VSS X110Y20VSSM VSS2 0.036nH
Rbump_X110Y30VDD X110Y30VDD X110Y30VDDM 20mOhm
Lbump_X110Y30VDD X110Y30VDDM VDD2 0.036nH
Rbump_X110Y30VSS X110Y30VSS X110Y30VSSM 20mOhm
Lbump_X110Y30VSS X110Y30VSSM VSS2 0.036nH
Rbump_X110Y40VDD X110Y40VDD X110Y40VDDM 20mOhm
Lbump_X110Y40VDD X110Y40VDDM VDD2 0.036nH
Rbump_X110Y40VSS X110Y40VSS X110Y40VSSM 20mOhm
Lbump_X110Y40VSS X110Y40VSSM VSS2 0.036nH
Rbump_X110Y50VDD X110Y50VDD X110Y50VDDM 20mOhm
Lbump_X110Y50VDD X110Y50VDDM VDD2 0.036nH
Rbump_X110Y50VSS X110Y50VSS X110Y50VSSM 20mOhm
Lbump_X110Y50VSS X110Y50VSSM VSS2 0.036nH
Rbump_X110Y60VDD X110Y60VDD X110Y60VDDM 20mOhm
Lbump_X110Y60VDD X110Y60VDDM VDD2 0.036nH
Rbump_X110Y60VSS X110Y60VSS X110Y60VSSM 20mOhm
Lbump_X110Y60VSS X110Y60VSSM VSS2 0.036nH
Rbump_X110Y70VDD X110Y70VDD X110Y70VDDM 20mOhm
Lbump_X110Y70VDD X110Y70VDDM VDD2 0.036nH
Rbump_X110Y70VSS X110Y70VSS X110Y70VSSM 20mOhm
Lbump_X110Y70VSS X110Y70VSSM VSS2 0.036nH
Rbump_X110Y80VDD X110Y80VDD X110Y80VDDM 20mOhm
Lbump_X110Y80VDD X110Y80VDDM VDD2 0.036nH
Rbump_X110Y80VSS X110Y80VSS X110Y80VSSM 20mOhm
Lbump_X110Y80VSS X110Y80VSSM VSS2 0.036nH
Rbump_X110Y90VDD X110Y90VDD X110Y90VDDM 20mOhm
Lbump_X110Y90VDD X110Y90VDDM VDD2 0.036nH
Rbump_X110Y90VSS X110Y90VSS X110Y90VSSM 20mOhm
Lbump_X110Y90VSS X110Y90VSSM VSS2 0.036nH
Rbump_X110Y100VDD X110Y100VDD X110Y100VDDM 20mOhm
Lbump_X110Y100VDD X110Y100VDDM VDD2 0.036nH
Rbump_X110Y100VSS X110Y100VSS X110Y100VSSM 20mOhm
Lbump_X110Y100VSS X110Y100VSSM VSS2 0.036nH
Rbump_X110Y110VDD X110Y110VDD X110Y110VDDM 20mOhm
Lbump_X110Y110VDD X110Y110VDDM VDD2 0.036nH
Rbump_X110Y110VSS X110Y110VSS X110Y110VSSM 20mOhm
Lbump_X110Y110VSS X110Y110VSSM VSS2 0.036nH
Rbump_X110Y120VDD X110Y120VDD X110Y120VDDM 20mOhm
Lbump_X110Y120VDD X110Y120VDDM VDD2 0.036nH
Rbump_X110Y120VSS X110Y120VSS X110Y120VSSM 20mOhm
Lbump_X110Y120VSS X110Y120VSSM VSS2 0.036nH
Rbump_X120Y10VDD X120Y10VDD X120Y10VDDM 20mOhm
Lbump_X120Y10VDD X120Y10VDDM VDD2 0.036nH
Rbump_X120Y10VSS X120Y10VSS X120Y10VSSM 20mOhm
Lbump_X120Y10VSS X120Y10VSSM VSS2 0.036nH
Rbump_X120Y20VDD X120Y20VDD X120Y20VDDM 20mOhm
Lbump_X120Y20VDD X120Y20VDDM VDD2 0.036nH
Rbump_X120Y20VSS X120Y20VSS X120Y20VSSM 20mOhm
Lbump_X120Y20VSS X120Y20VSSM VSS2 0.036nH
Rbump_X120Y30VDD X120Y30VDD X120Y30VDDM 20mOhm
Lbump_X120Y30VDD X120Y30VDDM VDD2 0.036nH
Rbump_X120Y30VSS X120Y30VSS X120Y30VSSM 20mOhm
Lbump_X120Y30VSS X120Y30VSSM VSS2 0.036nH
Rbump_X120Y40VDD X120Y40VDD X120Y40VDDM 20mOhm
Lbump_X120Y40VDD X120Y40VDDM VDD2 0.036nH
Rbump_X120Y40VSS X120Y40VSS X120Y40VSSM 20mOhm
Lbump_X120Y40VSS X120Y40VSSM VSS2 0.036nH
Rbump_X120Y50VDD X120Y50VDD X120Y50VDDM 20mOhm
Lbump_X120Y50VDD X120Y50VDDM VDD2 0.036nH
Rbump_X120Y50VSS X120Y50VSS X120Y50VSSM 20mOhm
Lbump_X120Y50VSS X120Y50VSSM VSS2 0.036nH
Rbump_X120Y60VDD X120Y60VDD X120Y60VDDM 20mOhm
Lbump_X120Y60VDD X120Y60VDDM VDD2 0.036nH
Rbump_X120Y60VSS X120Y60VSS X120Y60VSSM 20mOhm
Lbump_X120Y60VSS X120Y60VSSM VSS2 0.036nH
Rbump_X120Y70VDD X120Y70VDD X120Y70VDDM 20mOhm
Lbump_X120Y70VDD X120Y70VDDM VDD2 0.036nH
Rbump_X120Y70VSS X120Y70VSS X120Y70VSSM 20mOhm
Lbump_X120Y70VSS X120Y70VSSM VSS2 0.036nH
Rbump_X120Y80VDD X120Y80VDD X120Y80VDDM 20mOhm
Lbump_X120Y80VDD X120Y80VDDM VDD2 0.036nH
Rbump_X120Y80VSS X120Y80VSS X120Y80VSSM 20mOhm
Lbump_X120Y80VSS X120Y80VSSM VSS2 0.036nH
Rbump_X120Y90VDD X120Y90VDD X120Y90VDDM 20mOhm
Lbump_X120Y90VDD X120Y90VDDM VDD2 0.036nH
Rbump_X120Y90VSS X120Y90VSS X120Y90VSSM 20mOhm
Lbump_X120Y90VSS X120Y90VSSM VSS2 0.036nH
Rbump_X120Y100VDD X120Y100VDD X120Y100VDDM 20mOhm
Lbump_X120Y100VDD X120Y100VDDM VDD2 0.036nH
Rbump_X120Y100VSS X120Y100VSS X120Y100VSSM 20mOhm
Lbump_X120Y100VSS X120Y100VSSM VSS2 0.036nH
Rbump_X120Y110VDD X120Y110VDD X120Y110VDDM 20mOhm
Lbump_X120Y110VDD X120Y110VDDM VDD2 0.036nH
Rbump_X120Y110VSS X120Y110VSS X120Y110VSSM 20mOhm
Lbump_X120Y110VSS X120Y110VSSM VSS2 0.036nH
Rbump_X120Y120VDD X120Y120VDD X120Y120VDDM 20mOhm
Lbump_X120Y120VDD X120Y120VDDM VDD2 0.036nH
Rbump_X120Y120VSS X120Y120VSS X120Y120VSSM 20mOhm
Lbump_X120Y120VSS X120Y120VSSM VSS2 0.036nH
RsVDD VDD VDDMS 0.55mOhm
LsVDD VDDMS VDD2 0.06nH
RsVSS VSS VSSMS 0.55mOhm
LsVSS VSSMS VSS2 0.06nH
Rp VDD2 VDD2M 0.1mOhm
Lp VSS2 VSS2M 0.0028nH
Cp VDD2M VSS2M 52uF
.ends dut
XPcbBuckConverter0 VDD0 VSS0 PcbBuckConverter
Rgnd VSS0 0 0
XPcbModelLumped0 VDD0 VSS0 VDD1 VSS1 PcbModelLumped
Xdut VDD1 VSS1 dut


# case 1 distributed
.title 20200622-104933
.option rshunt = 1.0e12
.subckt Regulator VDD VSS
Vs VDD VSS 1.1
.ends Regulator

.subckt ChipPackage VDD1 VSS1 VDD2 VSS2
RsVDD VDD1 VDDMS 0.55mOhm
LsVDD VDDMS VDD2 0.06nH
RsVSS VSS1 VSSMS 0.55mOhm
LsVSS VSSMS VSS2 0.06nH
Rp VDD2 VDD2M 0.1mOhm
Lp VSS2 VSS2M 0.0028nH
Cp VDD2M VSS2M 52uF
.ends ChipPackage

.subckt ChipBump VDD1 VSS1 VDD2 VSS2
RX0Y0VDD VDD1 X0Y0VDDM 20mOhm
LX0Y0VDD X0Y0VDDM VDD2 0.036nH
RX0Y0VSS VSS1 X0Y0VSSM 20mOhm
LX0Y0VSS X0Y0VSSM VSS2 0.036nH
RX0Y1VDD VDD1 X0Y1VDDM 20mOhm
LX0Y1VDD X0Y1VDDM VDD2 0.036nH
RX0Y1VSS VSS1 X0Y1VSSM 20mOhm
LX0Y1VSS X0Y1VSSM VSS2 0.036nH
RX0Y2VDD VDD1 X0Y2VDDM 20mOhm
LX0Y2VDD X0Y2VDDM VDD2 0.036nH
RX0Y2VSS VSS1 X0Y2VSSM 20mOhm
LX0Y2VSS X0Y2VSSM VSS2 0.036nH
RX0Y3VDD VDD1 X0Y3VDDM 20mOhm
LX0Y3VDD X0Y3VDDM VDD2 0.036nH
RX0Y3VSS VSS1 X0Y3VSSM 20mOhm
LX0Y3VSS X0Y3VSSM VSS2 0.036nH
RX0Y4VDD VDD1 X0Y4VDDM 20mOhm
LX0Y4VDD X0Y4VDDM VDD2 0.036nH
RX0Y4VSS VSS1 X0Y4VSSM 20mOhm
LX0Y4VSS X0Y4VSSM VSS2 0.036nH
RX0Y5VDD VDD1 X0Y5VDDM 20mOhm
LX0Y5VDD X0Y5VDDM VDD2 0.036nH
RX0Y5VSS VSS1 X0Y5VSSM 20mOhm
LX0Y5VSS X0Y5VSSM VSS2 0.036nH
RX0Y6VDD VDD1 X0Y6VDDM 20mOhm
LX0Y6VDD X0Y6VDDM VDD2 0.036nH
RX0Y6VSS VSS1 X0Y6VSSM 20mOhm
LX0Y6VSS X0Y6VSSM VSS2 0.036nH
RX0Y7VDD VDD1 X0Y7VDDM 20mOhm
LX0Y7VDD X0Y7VDDM VDD2 0.036nH
RX0Y7VSS VSS1 X0Y7VSSM 20mOhm
LX0Y7VSS X0Y7VSSM VSS2 0.036nH
RX0Y8VDD VDD1 X0Y8VDDM 20mOhm
LX0Y8VDD X0Y8VDDM VDD2 0.036nH
RX0Y8VSS VSS1 X0Y8VSSM 20mOhm
LX0Y8VSS X0Y8VSSM VSS2 0.036nH
RX0Y9VDD VDD1 X0Y9VDDM 20mOhm
LX0Y9VDD X0Y9VDDM VDD2 0.036nH
RX0Y9VSS VSS1 X0Y9VSSM 20mOhm
LX0Y9VSS X0Y9VSSM VSS2 0.036nH
RX0Y10VDD VDD1 X0Y10VDDM 20mOhm
LX0Y10VDD X0Y10VDDM VDD2 0.036nH
RX0Y10VSS VSS1 X0Y10VSSM 20mOhm
LX0Y10VSS X0Y10VSSM VSS2 0.036nH
RX0Y11VDD VDD1 X0Y11VDDM 20mOhm
LX0Y11VDD X0Y11VDDM VDD2 0.036nH
RX0Y11VSS VSS1 X0Y11VSSM 20mOhm
LX0Y11VSS X0Y11VSSM VSS2 0.036nH
RX1Y0VDD VDD1 X1Y0VDDM 20mOhm
LX1Y0VDD X1Y0VDDM VDD2 0.036nH
RX1Y0VSS VSS1 X1Y0VSSM 20mOhm
LX1Y0VSS X1Y0VSSM VSS2 0.036nH
RX1Y1VDD VDD1 X1Y1VDDM 20mOhm
LX1Y1VDD X1Y1VDDM VDD2 0.036nH
RX1Y1VSS VSS1 X1Y1VSSM 20mOhm
LX1Y1VSS X1Y1VSSM VSS2 0.036nH
RX1Y2VDD VDD1 X1Y2VDDM 20mOhm
LX1Y2VDD X1Y2VDDM VDD2 0.036nH
RX1Y2VSS VSS1 X1Y2VSSM 20mOhm
LX1Y2VSS X1Y2VSSM VSS2 0.036nH
RX1Y3VDD VDD1 X1Y3VDDM 20mOhm
LX1Y3VDD X1Y3VDDM VDD2 0.036nH
RX1Y3VSS VSS1 X1Y3VSSM 20mOhm
LX1Y3VSS X1Y3VSSM VSS2 0.036nH
RX1Y4VDD VDD1 X1Y4VDDM 20mOhm
LX1Y4VDD X1Y4VDDM VDD2 0.036nH
RX1Y4VSS VSS1 X1Y4VSSM 20mOhm
LX1Y4VSS X1Y4VSSM VSS2 0.036nH
RX1Y5VDD VDD1 X1Y5VDDM 20mOhm
LX1Y5VDD X1Y5VDDM VDD2 0.036nH
RX1Y5VSS VSS1 X1Y5VSSM 20mOhm
LX1Y5VSS X1Y5VSSM VSS2 0.036nH
RX1Y6VDD VDD1 X1Y6VDDM 20mOhm
LX1Y6VDD X1Y6VDDM VDD2 0.036nH
RX1Y6VSS VSS1 X1Y6VSSM 20mOhm
LX1Y6VSS X1Y6VSSM VSS2 0.036nH
RX1Y7VDD VDD1 X1Y7VDDM 20mOhm
LX1Y7VDD X1Y7VDDM VDD2 0.036nH
RX1Y7VSS VSS1 X1Y7VSSM 20mOhm
LX1Y7VSS X1Y7VSSM VSS2 0.036nH
RX1Y8VDD VDD1 X1Y8VDDM 20mOhm
LX1Y8VDD X1Y8VDDM VDD2 0.036nH
RX1Y8VSS VSS1 X1Y8VSSM 20mOhm
LX1Y8VSS X1Y8VSSM VSS2 0.036nH
RX1Y9VDD VDD1 X1Y9VDDM 20mOhm
LX1Y9VDD X1Y9VDDM VDD2 0.036nH
RX1Y9VSS VSS1 X1Y9VSSM 20mOhm
LX1Y9VSS X1Y9VSSM VSS2 0.036nH
RX1Y10VDD VDD1 X1Y10VDDM 20mOhm
LX1Y10VDD X1Y10VDDM VDD2 0.036nH
RX1Y10VSS VSS1 X1Y10VSSM 20mOhm
LX1Y10VSS X1Y10VSSM VSS2 0.036nH
RX1Y11VDD VDD1 X1Y11VDDM 20mOhm
LX1Y11VDD X1Y11VDDM VDD2 0.036nH
RX1Y11VSS VSS1 X1Y11VSSM 20mOhm
LX1Y11VSS X1Y11VSSM VSS2 0.036nH
RX2Y0VDD VDD1 X2Y0VDDM 20mOhm
LX2Y0VDD X2Y0VDDM VDD2 0.036nH
RX2Y0VSS VSS1 X2Y0VSSM 20mOhm
LX2Y0VSS X2Y0VSSM VSS2 0.036nH
RX2Y1VDD VDD1 X2Y1VDDM 20mOhm
LX2Y1VDD X2Y1VDDM VDD2 0.036nH
RX2Y1VSS VSS1 X2Y1VSSM 20mOhm
LX2Y1VSS X2Y1VSSM VSS2 0.036nH
RX2Y2VDD VDD1 X2Y2VDDM 20mOhm
LX2Y2VDD X2Y2VDDM VDD2 0.036nH
RX2Y2VSS VSS1 X2Y2VSSM 20mOhm
LX2Y2VSS X2Y2VSSM VSS2 0.036nH
RX2Y3VDD VDD1 X2Y3VDDM 20mOhm
LX2Y3VDD X2Y3VDDM VDD2 0.036nH
RX2Y3VSS VSS1 X2Y3VSSM 20mOhm
LX2Y3VSS X2Y3VSSM VSS2 0.036nH
RX2Y4VDD VDD1 X2Y4VDDM 20mOhm
LX2Y4VDD X2Y4VDDM VDD2 0.036nH
RX2Y4VSS VSS1 X2Y4VSSM 20mOhm
LX2Y4VSS X2Y4VSSM VSS2 0.036nH
RX2Y5VDD VDD1 X2Y5VDDM 20mOhm
LX2Y5VDD X2Y5VDDM VDD2 0.036nH
RX2Y5VSS VSS1 X2Y5VSSM 20mOhm
LX2Y5VSS X2Y5VSSM VSS2 0.036nH
RX2Y6VDD VDD1 X2Y6VDDM 20mOhm
LX2Y6VDD X2Y6VDDM VDD2 0.036nH
RX2Y6VSS VSS1 X2Y6VSSM 20mOhm
LX2Y6VSS X2Y6VSSM VSS2 0.036nH
RX2Y7VDD VDD1 X2Y7VDDM 20mOhm
LX2Y7VDD X2Y7VDDM VDD2 0.036nH
RX2Y7VSS VSS1 X2Y7VSSM 20mOhm
LX2Y7VSS X2Y7VSSM VSS2 0.036nH
RX2Y8VDD VDD1 X2Y8VDDM 20mOhm
LX2Y8VDD X2Y8VDDM VDD2 0.036nH
RX2Y8VSS VSS1 X2Y8VSSM 20mOhm
LX2Y8VSS X2Y8VSSM VSS2 0.036nH
RX2Y9VDD VDD1 X2Y9VDDM 20mOhm
LX2Y9VDD X2Y9VDDM VDD2 0.036nH
RX2Y9VSS VSS1 X2Y9VSSM 20mOhm
LX2Y9VSS X2Y9VSSM VSS2 0.036nH
RX2Y10VDD VDD1 X2Y10VDDM 20mOhm
LX2Y10VDD X2Y10VDDM VDD2 0.036nH
RX2Y10VSS VSS1 X2Y10VSSM 20mOhm
LX2Y10VSS X2Y10VSSM VSS2 0.036nH
RX2Y11VDD VDD1 X2Y11VDDM 20mOhm
LX2Y11VDD X2Y11VDDM VDD2 0.036nH
RX2Y11VSS VSS1 X2Y11VSSM 20mOhm
LX2Y11VSS X2Y11VSSM VSS2 0.036nH
RX3Y0VDD VDD1 X3Y0VDDM 20mOhm
LX3Y0VDD X3Y0VDDM VDD2 0.036nH
RX3Y0VSS VSS1 X3Y0VSSM 20mOhm
LX3Y0VSS X3Y0VSSM VSS2 0.036nH
RX3Y1VDD VDD1 X3Y1VDDM 20mOhm
LX3Y1VDD X3Y1VDDM VDD2 0.036nH
RX3Y1VSS VSS1 X3Y1VSSM 20mOhm
LX3Y1VSS X3Y1VSSM VSS2 0.036nH
RX3Y2VDD VDD1 X3Y2VDDM 20mOhm
LX3Y2VDD X3Y2VDDM VDD2 0.036nH
RX3Y2VSS VSS1 X3Y2VSSM 20mOhm
LX3Y2VSS X3Y2VSSM VSS2 0.036nH
RX3Y3VDD VDD1 X3Y3VDDM 20mOhm
LX3Y3VDD X3Y3VDDM VDD2 0.036nH
RX3Y3VSS VSS1 X3Y3VSSM 20mOhm
LX3Y3VSS X3Y3VSSM VSS2 0.036nH
RX3Y4VDD VDD1 X3Y4VDDM 20mOhm
LX3Y4VDD X3Y4VDDM VDD2 0.036nH
RX3Y4VSS VSS1 X3Y4VSSM 20mOhm
LX3Y4VSS X3Y4VSSM VSS2 0.036nH
RX3Y5VDD VDD1 X3Y5VDDM 20mOhm
LX3Y5VDD X3Y5VDDM VDD2 0.036nH
RX3Y5VSS VSS1 X3Y5VSSM 20mOhm
LX3Y5VSS X3Y5VSSM VSS2 0.036nH
RX3Y6VDD VDD1 X3Y6VDDM 20mOhm
LX3Y6VDD X3Y6VDDM VDD2 0.036nH
RX3Y6VSS VSS1 X3Y6VSSM 20mOhm
LX3Y6VSS X3Y6VSSM VSS2 0.036nH
RX3Y7VDD VDD1 X3Y7VDDM 20mOhm
LX3Y7VDD X3Y7VDDM VDD2 0.036nH
RX3Y7VSS VSS1 X3Y7VSSM 20mOhm
LX3Y7VSS X3Y7VSSM VSS2 0.036nH
RX3Y8VDD VDD1 X3Y8VDDM 20mOhm
LX3Y8VDD X3Y8VDDM VDD2 0.036nH
RX3Y8VSS VSS1 X3Y8VSSM 20mOhm
LX3Y8VSS X3Y8VSSM VSS2 0.036nH
RX3Y9VDD VDD1 X3Y9VDDM 20mOhm
LX3Y9VDD X3Y9VDDM VDD2 0.036nH
RX3Y9VSS VSS1 X3Y9VSSM 20mOhm
LX3Y9VSS X3Y9VSSM VSS2 0.036nH
RX3Y10VDD VDD1 X3Y10VDDM 20mOhm
LX3Y10VDD X3Y10VDDM VDD2 0.036nH
RX3Y10VSS VSS1 X3Y10VSSM 20mOhm
LX3Y10VSS X3Y10VSSM VSS2 0.036nH
RX3Y11VDD VDD1 X3Y11VDDM 20mOhm
LX3Y11VDD X3Y11VDDM VDD2 0.036nH
RX3Y11VSS VSS1 X3Y11VSSM 20mOhm
LX3Y11VSS X3Y11VSSM VSS2 0.036nH
RX4Y0VDD VDD1 X4Y0VDDM 20mOhm
LX4Y0VDD X4Y0VDDM VDD2 0.036nH
RX4Y0VSS VSS1 X4Y0VSSM 20mOhm
LX4Y0VSS X4Y0VSSM VSS2 0.036nH
RX4Y1VDD VDD1 X4Y1VDDM 20mOhm
LX4Y1VDD X4Y1VDDM VDD2 0.036nH
RX4Y1VSS VSS1 X4Y1VSSM 20mOhm
LX4Y1VSS X4Y1VSSM VSS2 0.036nH
RX4Y2VDD VDD1 X4Y2VDDM 20mOhm
LX4Y2VDD X4Y2VDDM VDD2 0.036nH
RX4Y2VSS VSS1 X4Y2VSSM 20mOhm
LX4Y2VSS X4Y2VSSM VSS2 0.036nH
RX4Y3VDD VDD1 X4Y3VDDM 20mOhm
LX4Y3VDD X4Y3VDDM VDD2 0.036nH
RX4Y3VSS VSS1 X4Y3VSSM 20mOhm
LX4Y3VSS X4Y3VSSM VSS2 0.036nH
RX4Y4VDD VDD1 X4Y4VDDM 20mOhm
LX4Y4VDD X4Y4VDDM VDD2 0.036nH
RX4Y4VSS VSS1 X4Y4VSSM 20mOhm
LX4Y4VSS X4Y4VSSM VSS2 0.036nH
RX4Y5VDD VDD1 X4Y5VDDM 20mOhm
LX4Y5VDD X4Y5VDDM VDD2 0.036nH
RX4Y5VSS VSS1 X4Y5VSSM 20mOhm
LX4Y5VSS X4Y5VSSM VSS2 0.036nH
RX4Y6VDD VDD1 X4Y6VDDM 20mOhm
LX4Y6VDD X4Y6VDDM VDD2 0.036nH
RX4Y6VSS VSS1 X4Y6VSSM 20mOhm
LX4Y6VSS X4Y6VSSM VSS2 0.036nH
RX4Y7VDD VDD1 X4Y7VDDM 20mOhm
LX4Y7VDD X4Y7VDDM VDD2 0.036nH
RX4Y7VSS VSS1 X4Y7VSSM 20mOhm
LX4Y7VSS X4Y7VSSM VSS2 0.036nH
RX4Y8VDD VDD1 X4Y8VDDM 20mOhm
LX4Y8VDD X4Y8VDDM VDD2 0.036nH
RX4Y8VSS VSS1 X4Y8VSSM 20mOhm
LX4Y8VSS X4Y8VSSM VSS2 0.036nH
RX4Y9VDD VDD1 X4Y9VDDM 20mOhm
LX4Y9VDD X4Y9VDDM VDD2 0.036nH
RX4Y9VSS VSS1 X4Y9VSSM 20mOhm
LX4Y9VSS X4Y9VSSM VSS2 0.036nH
RX4Y10VDD VDD1 X4Y10VDDM 20mOhm
LX4Y10VDD X4Y10VDDM VDD2 0.036nH
RX4Y10VSS VSS1 X4Y10VSSM 20mOhm
LX4Y10VSS X4Y10VSSM VSS2 0.036nH
RX4Y11VDD VDD1 X4Y11VDDM 20mOhm
LX4Y11VDD X4Y11VDDM VDD2 0.036nH
RX4Y11VSS VSS1 X4Y11VSSM 20mOhm
LX4Y11VSS X4Y11VSSM VSS2 0.036nH
RX5Y0VDD VDD1 X5Y0VDDM 20mOhm
LX5Y0VDD X5Y0VDDM VDD2 0.036nH
RX5Y0VSS VSS1 X5Y0VSSM 20mOhm
LX5Y0VSS X5Y0VSSM VSS2 0.036nH
RX5Y1VDD VDD1 X5Y1VDDM 20mOhm
LX5Y1VDD X5Y1VDDM VDD2 0.036nH
RX5Y1VSS VSS1 X5Y1VSSM 20mOhm
LX5Y1VSS X5Y1VSSM VSS2 0.036nH
RX5Y2VDD VDD1 X5Y2VDDM 20mOhm
LX5Y2VDD X5Y2VDDM VDD2 0.036nH
RX5Y2VSS VSS1 X5Y2VSSM 20mOhm
LX5Y2VSS X5Y2VSSM VSS2 0.036nH
RX5Y3VDD VDD1 X5Y3VDDM 20mOhm
LX5Y3VDD X5Y3VDDM VDD2 0.036nH
RX5Y3VSS VSS1 X5Y3VSSM 20mOhm
LX5Y3VSS X5Y3VSSM VSS2 0.036nH
RX5Y4VDD VDD1 X5Y4VDDM 20mOhm
LX5Y4VDD X5Y4VDDM VDD2 0.036nH
RX5Y4VSS VSS1 X5Y4VSSM 20mOhm
LX5Y4VSS X5Y4VSSM VSS2 0.036nH
RX5Y5VDD VDD1 X5Y5VDDM 20mOhm
LX5Y5VDD X5Y5VDDM VDD2 0.036nH
RX5Y5VSS VSS1 X5Y5VSSM 20mOhm
LX5Y5VSS X5Y5VSSM VSS2 0.036nH
RX5Y6VDD VDD1 X5Y6VDDM 20mOhm
LX5Y6VDD X5Y6VDDM VDD2 0.036nH
RX5Y6VSS VSS1 X5Y6VSSM 20mOhm
LX5Y6VSS X5Y6VSSM VSS2 0.036nH
RX5Y7VDD VDD1 X5Y7VDDM 20mOhm
LX5Y7VDD X5Y7VDDM VDD2 0.036nH
RX5Y7VSS VSS1 X5Y7VSSM 20mOhm
LX5Y7VSS X5Y7VSSM VSS2 0.036nH
RX5Y8VDD VDD1 X5Y8VDDM 20mOhm
LX5Y8VDD X5Y8VDDM VDD2 0.036nH
RX5Y8VSS VSS1 X5Y8VSSM 20mOhm
LX5Y8VSS X5Y8VSSM VSS2 0.036nH
RX5Y9VDD VDD1 X5Y9VDDM 20mOhm
LX5Y9VDD X5Y9VDDM VDD2 0.036nH
RX5Y9VSS VSS1 X5Y9VSSM 20mOhm
LX5Y9VSS X5Y9VSSM VSS2 0.036nH
RX5Y10VDD VDD1 X5Y10VDDM 20mOhm
LX5Y10VDD X5Y10VDDM VDD2 0.036nH
RX5Y10VSS VSS1 X5Y10VSSM 20mOhm
LX5Y10VSS X5Y10VSSM VSS2 0.036nH
RX5Y11VDD VDD1 X5Y11VDDM 20mOhm
LX5Y11VDD X5Y11VDDM VDD2 0.036nH
RX5Y11VSS VSS1 X5Y11VSSM 20mOhm
LX5Y11VSS X5Y11VSSM VSS2 0.036nH
RX6Y0VDD VDD1 X6Y0VDDM 20mOhm
LX6Y0VDD X6Y0VDDM VDD2 0.036nH
RX6Y0VSS VSS1 X6Y0VSSM 20mOhm
LX6Y0VSS X6Y0VSSM VSS2 0.036nH
RX6Y1VDD VDD1 X6Y1VDDM 20mOhm
LX6Y1VDD X6Y1VDDM VDD2 0.036nH
RX6Y1VSS VSS1 X6Y1VSSM 20mOhm
LX6Y1VSS X6Y1VSSM VSS2 0.036nH
RX6Y2VDD VDD1 X6Y2VDDM 20mOhm
LX6Y2VDD X6Y2VDDM VDD2 0.036nH
RX6Y2VSS VSS1 X6Y2VSSM 20mOhm
LX6Y2VSS X6Y2VSSM VSS2 0.036nH
RX6Y3VDD VDD1 X6Y3VDDM 20mOhm
LX6Y3VDD X6Y3VDDM VDD2 0.036nH
RX6Y3VSS VSS1 X6Y3VSSM 20mOhm
LX6Y3VSS X6Y3VSSM VSS2 0.036nH
RX6Y4VDD VDD1 X6Y4VDDM 20mOhm
LX6Y4VDD X6Y4VDDM VDD2 0.036nH
RX6Y4VSS VSS1 X6Y4VSSM 20mOhm
LX6Y4VSS X6Y4VSSM VSS2 0.036nH
RX6Y5VDD VDD1 X6Y5VDDM 20mOhm
LX6Y5VDD X6Y5VDDM VDD2 0.036nH
RX6Y5VSS VSS1 X6Y5VSSM 20mOhm
LX6Y5VSS X6Y5VSSM VSS2 0.036nH
RX6Y6VDD VDD1 X6Y6VDDM 20mOhm
LX6Y6VDD X6Y6VDDM VDD2 0.036nH
RX6Y6VSS VSS1 X6Y6VSSM 20mOhm
LX6Y6VSS X6Y6VSSM VSS2 0.036nH
RX6Y7VDD VDD1 X6Y7VDDM 20mOhm
LX6Y7VDD X6Y7VDDM VDD2 0.036nH
RX6Y7VSS VSS1 X6Y7VSSM 20mOhm
LX6Y7VSS X6Y7VSSM VSS2 0.036nH
RX6Y8VDD VDD1 X6Y8VDDM 20mOhm
LX6Y8VDD X6Y8VDDM VDD2 0.036nH
RX6Y8VSS VSS1 X6Y8VSSM 20mOhm
LX6Y8VSS X6Y8VSSM VSS2 0.036nH
RX6Y9VDD VDD1 X6Y9VDDM 20mOhm
LX6Y9VDD X6Y9VDDM VDD2 0.036nH
RX6Y9VSS VSS1 X6Y9VSSM 20mOhm
LX6Y9VSS X6Y9VSSM VSS2 0.036nH
RX6Y10VDD VDD1 X6Y10VDDM 20mOhm
LX6Y10VDD X6Y10VDDM VDD2 0.036nH
RX6Y10VSS VSS1 X6Y10VSSM 20mOhm
LX6Y10VSS X6Y10VSSM VSS2 0.036nH
RX6Y11VDD VDD1 X6Y11VDDM 20mOhm
LX6Y11VDD X6Y11VDDM VDD2 0.036nH
RX6Y11VSS VSS1 X6Y11VSSM 20mOhm
LX6Y11VSS X6Y11VSSM VSS2 0.036nH
RX7Y0VDD VDD1 X7Y0VDDM 20mOhm
LX7Y0VDD X7Y0VDDM VDD2 0.036nH
RX7Y0VSS VSS1 X7Y0VSSM 20mOhm
LX7Y0VSS X7Y0VSSM VSS2 0.036nH
RX7Y1VDD VDD1 X7Y1VDDM 20mOhm
LX7Y1VDD X7Y1VDDM VDD2 0.036nH
RX7Y1VSS VSS1 X7Y1VSSM 20mOhm
LX7Y1VSS X7Y1VSSM VSS2 0.036nH
RX7Y2VDD VDD1 X7Y2VDDM 20mOhm
LX7Y2VDD X7Y2VDDM VDD2 0.036nH
RX7Y2VSS VSS1 X7Y2VSSM 20mOhm
LX7Y2VSS X7Y2VSSM VSS2 0.036nH
RX7Y3VDD VDD1 X7Y3VDDM 20mOhm
LX7Y3VDD X7Y3VDDM VDD2 0.036nH
RX7Y3VSS VSS1 X7Y3VSSM 20mOhm
LX7Y3VSS X7Y3VSSM VSS2 0.036nH
RX7Y4VDD VDD1 X7Y4VDDM 20mOhm
LX7Y4VDD X7Y4VDDM VDD2 0.036nH
RX7Y4VSS VSS1 X7Y4VSSM 20mOhm
LX7Y4VSS X7Y4VSSM VSS2 0.036nH
RX7Y5VDD VDD1 X7Y5VDDM 20mOhm
LX7Y5VDD X7Y5VDDM VDD2 0.036nH
RX7Y5VSS VSS1 X7Y5VSSM 20mOhm
LX7Y5VSS X7Y5VSSM VSS2 0.036nH
RX7Y6VDD VDD1 X7Y6VDDM 20mOhm
LX7Y6VDD X7Y6VDDM VDD2 0.036nH
RX7Y6VSS VSS1 X7Y6VSSM 20mOhm
LX7Y6VSS X7Y6VSSM VSS2 0.036nH
RX7Y7VDD VDD1 X7Y7VDDM 20mOhm
LX7Y7VDD X7Y7VDDM VDD2 0.036nH
RX7Y7VSS VSS1 X7Y7VSSM 20mOhm
LX7Y7VSS X7Y7VSSM VSS2 0.036nH
RX7Y8VDD VDD1 X7Y8VDDM 20mOhm
LX7Y8VDD X7Y8VDDM VDD2 0.036nH
RX7Y8VSS VSS1 X7Y8VSSM 20mOhm
LX7Y8VSS X7Y8VSSM VSS2 0.036nH
RX7Y9VDD VDD1 X7Y9VDDM 20mOhm
LX7Y9VDD X7Y9VDDM VDD2 0.036nH
RX7Y9VSS VSS1 X7Y9VSSM 20mOhm
LX7Y9VSS X7Y9VSSM VSS2 0.036nH
RX7Y10VDD VDD1 X7Y10VDDM 20mOhm
LX7Y10VDD X7Y10VDDM VDD2 0.036nH
RX7Y10VSS VSS1 X7Y10VSSM 20mOhm
LX7Y10VSS X7Y10VSSM VSS2 0.036nH
RX7Y11VDD VDD1 X7Y11VDDM 20mOhm
LX7Y11VDD X7Y11VDDM VDD2 0.036nH
RX7Y11VSS VSS1 X7Y11VSSM 20mOhm
LX7Y11VSS X7Y11VSSM VSS2 0.036nH
RX8Y0VDD VDD1 X8Y0VDDM 20mOhm
LX8Y0VDD X8Y0VDDM VDD2 0.036nH
RX8Y0VSS VSS1 X8Y0VSSM 20mOhm
LX8Y0VSS X8Y0VSSM VSS2 0.036nH
RX8Y1VDD VDD1 X8Y1VDDM 20mOhm
LX8Y1VDD X8Y1VDDM VDD2 0.036nH
RX8Y1VSS VSS1 X8Y1VSSM 20mOhm
LX8Y1VSS X8Y1VSSM VSS2 0.036nH
RX8Y2VDD VDD1 X8Y2VDDM 20mOhm
LX8Y2VDD X8Y2VDDM VDD2 0.036nH
RX8Y2VSS VSS1 X8Y2VSSM 20mOhm
LX8Y2VSS X8Y2VSSM VSS2 0.036nH
RX8Y3VDD VDD1 X8Y3VDDM 20mOhm
LX8Y3VDD X8Y3VDDM VDD2 0.036nH
RX8Y3VSS VSS1 X8Y3VSSM 20mOhm
LX8Y3VSS X8Y3VSSM VSS2 0.036nH
RX8Y4VDD VDD1 X8Y4VDDM 20mOhm
LX8Y4VDD X8Y4VDDM VDD2 0.036nH
RX8Y4VSS VSS1 X8Y4VSSM 20mOhm
LX8Y4VSS X8Y4VSSM VSS2 0.036nH
RX8Y5VDD VDD1 X8Y5VDDM 20mOhm
LX8Y5VDD X8Y5VDDM VDD2 0.036nH
RX8Y5VSS VSS1 X8Y5VSSM 20mOhm
LX8Y5VSS X8Y5VSSM VSS2 0.036nH
RX8Y6VDD VDD1 X8Y6VDDM 20mOhm
LX8Y6VDD X8Y6VDDM VDD2 0.036nH
RX8Y6VSS VSS1 X8Y6VSSM 20mOhm
LX8Y6VSS X8Y6VSSM VSS2 0.036nH
RX8Y7VDD VDD1 X8Y7VDDM 20mOhm
LX8Y7VDD X8Y7VDDM VDD2 0.036nH
RX8Y7VSS VSS1 X8Y7VSSM 20mOhm
LX8Y7VSS X8Y7VSSM VSS2 0.036nH
RX8Y8VDD VDD1 X8Y8VDDM 20mOhm
LX8Y8VDD X8Y8VDDM VDD2 0.036nH
RX8Y8VSS VSS1 X8Y8VSSM 20mOhm
LX8Y8VSS X8Y8VSSM VSS2 0.036nH
RX8Y9VDD VDD1 X8Y9VDDM 20mOhm
LX8Y9VDD X8Y9VDDM VDD2 0.036nH
RX8Y9VSS VSS1 X8Y9VSSM 20mOhm
LX8Y9VSS X8Y9VSSM VSS2 0.036nH
RX8Y10VDD VDD1 X8Y10VDDM 20mOhm
LX8Y10VDD X8Y10VDDM VDD2 0.036nH
RX8Y10VSS VSS1 X8Y10VSSM 20mOhm
LX8Y10VSS X8Y10VSSM VSS2 0.036nH
RX8Y11VDD VDD1 X8Y11VDDM 20mOhm
LX8Y11VDD X8Y11VDDM VDD2 0.036nH
RX8Y11VSS VSS1 X8Y11VSSM 20mOhm
LX8Y11VSS X8Y11VSSM VSS2 0.036nH
RX9Y0VDD VDD1 X9Y0VDDM 20mOhm
LX9Y0VDD X9Y0VDDM VDD2 0.036nH
RX9Y0VSS VSS1 X9Y0VSSM 20mOhm
LX9Y0VSS X9Y0VSSM VSS2 0.036nH
RX9Y1VDD VDD1 X9Y1VDDM 20mOhm
LX9Y1VDD X9Y1VDDM VDD2 0.036nH
RX9Y1VSS VSS1 X9Y1VSSM 20mOhm
LX9Y1VSS X9Y1VSSM VSS2 0.036nH
RX9Y2VDD VDD1 X9Y2VDDM 20mOhm
LX9Y2VDD X9Y2VDDM VDD2 0.036nH
RX9Y2VSS VSS1 X9Y2VSSM 20mOhm
LX9Y2VSS X9Y2VSSM VSS2 0.036nH
RX9Y3VDD VDD1 X9Y3VDDM 20mOhm
LX9Y3VDD X9Y3VDDM VDD2 0.036nH
RX9Y3VSS VSS1 X9Y3VSSM 20mOhm
LX9Y3VSS X9Y3VSSM VSS2 0.036nH
RX9Y4VDD VDD1 X9Y4VDDM 20mOhm
LX9Y4VDD X9Y4VDDM VDD2 0.036nH
RX9Y4VSS VSS1 X9Y4VSSM 20mOhm
LX9Y4VSS X9Y4VSSM VSS2 0.036nH
RX9Y5VDD VDD1 X9Y5VDDM 20mOhm
LX9Y5VDD X9Y5VDDM VDD2 0.036nH
RX9Y5VSS VSS1 X9Y5VSSM 20mOhm
LX9Y5VSS X9Y5VSSM VSS2 0.036nH
RX9Y6VDD VDD1 X9Y6VDDM 20mOhm
LX9Y6VDD X9Y6VDDM VDD2 0.036nH
RX9Y6VSS VSS1 X9Y6VSSM 20mOhm
LX9Y6VSS X9Y6VSSM VSS2 0.036nH
RX9Y7VDD VDD1 X9Y7VDDM 20mOhm
LX9Y7VDD X9Y7VDDM VDD2 0.036nH
RX9Y7VSS VSS1 X9Y7VSSM 20mOhm
LX9Y7VSS X9Y7VSSM VSS2 0.036nH
RX9Y8VDD VDD1 X9Y8VDDM 20mOhm
LX9Y8VDD X9Y8VDDM VDD2 0.036nH
RX9Y8VSS VSS1 X9Y8VSSM 20mOhm
LX9Y8VSS X9Y8VSSM VSS2 0.036nH
RX9Y9VDD VDD1 X9Y9VDDM 20mOhm
LX9Y9VDD X9Y9VDDM VDD2 0.036nH
RX9Y9VSS VSS1 X9Y9VSSM 20mOhm
LX9Y9VSS X9Y9VSSM VSS2 0.036nH
RX9Y10VDD VDD1 X9Y10VDDM 20mOhm
LX9Y10VDD X9Y10VDDM VDD2 0.036nH
RX9Y10VSS VSS1 X9Y10VSSM 20mOhm
LX9Y10VSS X9Y10VSSM VSS2 0.036nH
RX9Y11VDD VDD1 X9Y11VDDM 20mOhm
LX9Y11VDD X9Y11VDDM VDD2 0.036nH
RX9Y11VSS VSS1 X9Y11VSSM 20mOhm
LX9Y11VSS X9Y11VSSM VSS2 0.036nH
RX10Y0VDD VDD1 X10Y0VDDM 20mOhm
LX10Y0VDD X10Y0VDDM VDD2 0.036nH
RX10Y0VSS VSS1 X10Y0VSSM 20mOhm
LX10Y0VSS X10Y0VSSM VSS2 0.036nH
RX10Y1VDD VDD1 X10Y1VDDM 20mOhm
LX10Y1VDD X10Y1VDDM VDD2 0.036nH
RX10Y1VSS VSS1 X10Y1VSSM 20mOhm
LX10Y1VSS X10Y1VSSM VSS2 0.036nH
RX10Y2VDD VDD1 X10Y2VDDM 20mOhm
LX10Y2VDD X10Y2VDDM VDD2 0.036nH
RX10Y2VSS VSS1 X10Y2VSSM 20mOhm
LX10Y2VSS X10Y2VSSM VSS2 0.036nH
RX10Y3VDD VDD1 X10Y3VDDM 20mOhm
LX10Y3VDD X10Y3VDDM VDD2 0.036nH
RX10Y3VSS VSS1 X10Y3VSSM 20mOhm
LX10Y3VSS X10Y3VSSM VSS2 0.036nH
RX10Y4VDD VDD1 X10Y4VDDM 20mOhm
LX10Y4VDD X10Y4VDDM VDD2 0.036nH
RX10Y4VSS VSS1 X10Y4VSSM 20mOhm
LX10Y4VSS X10Y4VSSM VSS2 0.036nH
RX10Y5VDD VDD1 X10Y5VDDM 20mOhm
LX10Y5VDD X10Y5VDDM VDD2 0.036nH
RX10Y5VSS VSS1 X10Y5VSSM 20mOhm
LX10Y5VSS X10Y5VSSM VSS2 0.036nH
RX10Y6VDD VDD1 X10Y6VDDM 20mOhm
LX10Y6VDD X10Y6VDDM VDD2 0.036nH
RX10Y6VSS VSS1 X10Y6VSSM 20mOhm
LX10Y6VSS X10Y6VSSM VSS2 0.036nH
RX10Y7VDD VDD1 X10Y7VDDM 20mOhm
LX10Y7VDD X10Y7VDDM VDD2 0.036nH
RX10Y7VSS VSS1 X10Y7VSSM 20mOhm
LX10Y7VSS X10Y7VSSM VSS2 0.036nH
RX10Y8VDD VDD1 X10Y8VDDM 20mOhm
LX10Y8VDD X10Y8VDDM VDD2 0.036nH
RX10Y8VSS VSS1 X10Y8VSSM 20mOhm
LX10Y8VSS X10Y8VSSM VSS2 0.036nH
RX10Y9VDD VDD1 X10Y9VDDM 20mOhm
LX10Y9VDD X10Y9VDDM VDD2 0.036nH
RX10Y9VSS VSS1 X10Y9VSSM 20mOhm
LX10Y9VSS X10Y9VSSM VSS2 0.036nH
RX10Y10VDD VDD1 X10Y10VDDM 20mOhm
LX10Y10VDD X10Y10VDDM VDD2 0.036nH
RX10Y10VSS VSS1 X10Y10VSSM 20mOhm
LX10Y10VSS X10Y10VSSM VSS2 0.036nH
RX10Y11VDD VDD1 X10Y11VDDM 20mOhm
LX10Y11VDD X10Y11VDDM VDD2 0.036nH
RX10Y11VSS VSS1 X10Y11VSSM 20mOhm
LX10Y11VSS X10Y11VSSM VSS2 0.036nH
RX11Y0VDD VDD1 X11Y0VDDM 20mOhm
LX11Y0VDD X11Y0VDDM VDD2 0.036nH
RX11Y0VSS VSS1 X11Y0VSSM 20mOhm
LX11Y0VSS X11Y0VSSM VSS2 0.036nH
RX11Y1VDD VDD1 X11Y1VDDM 20mOhm
LX11Y1VDD X11Y1VDDM VDD2 0.036nH
RX11Y1VSS VSS1 X11Y1VSSM 20mOhm
LX11Y1VSS X11Y1VSSM VSS2 0.036nH
RX11Y2VDD VDD1 X11Y2VDDM 20mOhm
LX11Y2VDD X11Y2VDDM VDD2 0.036nH
RX11Y2VSS VSS1 X11Y2VSSM 20mOhm
LX11Y2VSS X11Y2VSSM VSS2 0.036nH
RX11Y3VDD VDD1 X11Y3VDDM 20mOhm
LX11Y3VDD X11Y3VDDM VDD2 0.036nH
RX11Y3VSS VSS1 X11Y3VSSM 20mOhm
LX11Y3VSS X11Y3VSSM VSS2 0.036nH
RX11Y4VDD VDD1 X11Y4VDDM 20mOhm
LX11Y4VDD X11Y4VDDM VDD2 0.036nH
RX11Y4VSS VSS1 X11Y4VSSM 20mOhm
LX11Y4VSS X11Y4VSSM VSS2 0.036nH
RX11Y5VDD VDD1 X11Y5VDDM 20mOhm
LX11Y5VDD X11Y5VDDM VDD2 0.036nH
RX11Y5VSS VSS1 X11Y5VSSM 20mOhm
LX11Y5VSS X11Y5VSSM VSS2 0.036nH
RX11Y6VDD VDD1 X11Y6VDDM 20mOhm
LX11Y6VDD X11Y6VDDM VDD2 0.036nH
RX11Y6VSS VSS1 X11Y6VSSM 20mOhm
LX11Y6VSS X11Y6VSSM VSS2 0.036nH
RX11Y7VDD VDD1 X11Y7VDDM 20mOhm
LX11Y7VDD X11Y7VDDM VDD2 0.036nH
RX11Y7VSS VSS1 X11Y7VSSM 20mOhm
LX11Y7VSS X11Y7VSSM VSS2 0.036nH
RX11Y8VDD VDD1 X11Y8VDDM 20mOhm
LX11Y8VDD X11Y8VDDM VDD2 0.036nH
RX11Y8VSS VSS1 X11Y8VSSM 20mOhm
LX11Y8VSS X11Y8VSSM VSS2 0.036nH
RX11Y9VDD VDD1 X11Y9VDDM 20mOhm
LX11Y9VDD X11Y9VDDM VDD2 0.036nH
RX11Y9VSS VSS1 X11Y9VSSM 20mOhm
LX11Y9VSS X11Y9VSSM VSS2 0.036nH
RX11Y10VDD VDD1 X11Y10VDDM 20mOhm
LX11Y10VDD X11Y10VDDM VDD2 0.036nH
RX11Y10VSS VSS1 X11Y10VSSM 20mOhm
LX11Y10VSS X11Y10VSSM VSS2 0.036nH
RX11Y11VDD VDD1 X11Y11VDDM 20mOhm
LX11Y11VDD X11Y11VDDM VDD2 0.036nH
RX11Y11VSS VSS1 X11Y11VSSM 20mOhm
LX11Y11VSS X11Y11VSSM VSS2 0.036nH
.ends ChipBump

.subckt PcbModelLumped VDD1 VSS1 VDD2 VSS2
Rs1 VDD1 11 1000mOhm
Ls1 11 VDD2 0nH
Rs2 VSS1 21 1000mOhm
Ls2 21 VSS2 0nH
Rp VDD2 VDD2M 0mOhm
Cp VDD2M VSS2 0uF
.ends PcbModelLumped

.subckt dut VDD VSS
R_X10Y10VDD_X20Y10VDD X10Y10VDD X15Y10VDD 25mOhm
L_X10Y10VDD_X20Y10VDD X15Y10VDD X20Y10VDD 2.91e-06nH
R_X10Y10VSS_X20Y10VSS X10Y10VSS X15Y10VSS 25mOhm
L_X10Y10VSS_X20Y10VSS X15Y10VSS X20Y10VSS 2.91e-06nH
R_X20Y10VDD_X30Y10VDD X20Y10VDD X25Y10VDD 25mOhm
L_X20Y10VDD_X30Y10VDD X25Y10VDD X30Y10VDD 2.91e-06nH
R_X20Y10VSS_X30Y10VSS X20Y10VSS X25Y10VSS 25mOhm
L_X20Y10VSS_X30Y10VSS X25Y10VSS X30Y10VSS 2.91e-06nH
R_X30Y10VDD_X40Y10VDD X30Y10VDD X35Y10VDD 25mOhm
L_X30Y10VDD_X40Y10VDD X35Y10VDD X40Y10VDD 2.91e-06nH
R_X30Y10VSS_X40Y10VSS X30Y10VSS X35Y10VSS 25mOhm
L_X30Y10VSS_X40Y10VSS X35Y10VSS X40Y10VSS 2.91e-06nH
R_X40Y10VDD_X50Y10VDD X40Y10VDD X45Y10VDD 25mOhm
L_X40Y10VDD_X50Y10VDD X45Y10VDD X50Y10VDD 2.91e-06nH
R_X40Y10VSS_X50Y10VSS X40Y10VSS X45Y10VSS 25mOhm
L_X40Y10VSS_X50Y10VSS X45Y10VSS X50Y10VSS 2.91e-06nH
R_X50Y10VDD_X60Y10VDD X50Y10VDD X55Y10VDD 25mOhm
L_X50Y10VDD_X60Y10VDD X55Y10VDD X60Y10VDD 2.91e-06nH
R_X50Y10VSS_X60Y10VSS X50Y10VSS X55Y10VSS 25mOhm
L_X50Y10VSS_X60Y10VSS X55Y10VSS X60Y10VSS 2.91e-06nH
R_X60Y10VDD_X70Y10VDD X60Y10VDD X65Y10VDD 25mOhm
L_X60Y10VDD_X70Y10VDD X65Y10VDD X70Y10VDD 2.91e-06nH
R_X60Y10VSS_X70Y10VSS X60Y10VSS X65Y10VSS 25mOhm
L_X60Y10VSS_X70Y10VSS X65Y10VSS X70Y10VSS 2.91e-06nH
R_X70Y10VDD_X80Y10VDD X70Y10VDD X75Y10VDD 25mOhm
L_X70Y10VDD_X80Y10VDD X75Y10VDD X80Y10VDD 2.91e-06nH
R_X70Y10VSS_X80Y10VSS X70Y10VSS X75Y10VSS 25mOhm
L_X70Y10VSS_X80Y10VSS X75Y10VSS X80Y10VSS 2.91e-06nH
R_X80Y10VDD_X90Y10VDD X80Y10VDD X85Y10VDD 25mOhm
L_X80Y10VDD_X90Y10VDD X85Y10VDD X90Y10VDD 2.91e-06nH
R_X80Y10VSS_X90Y10VSS X80Y10VSS X85Y10VSS 25mOhm
L_X80Y10VSS_X90Y10VSS X85Y10VSS X90Y10VSS 2.91e-06nH
R_X90Y10VDD_X100Y10VDD X90Y10VDD X95Y10VDD 25mOhm
L_X90Y10VDD_X100Y10VDD X95Y10VDD X100Y10VDD 2.91e-06nH
R_X90Y10VSS_X100Y10VSS X90Y10VSS X95Y10VSS 25mOhm
L_X90Y10VSS_X100Y10VSS X95Y10VSS X100Y10VSS 2.91e-06nH
R_X100Y10VDD_X110Y10VDD X100Y10VDD X105Y10VDD 25mOhm
L_X100Y10VDD_X110Y10VDD X105Y10VDD X110Y10VDD 2.91e-06nH
R_X100Y10VSS_X110Y10VSS X100Y10VSS X105Y10VSS 25mOhm
L_X100Y10VSS_X110Y10VSS X105Y10VSS X110Y10VSS 2.91e-06nH
R_X110Y10VDD_X120Y10VDD X110Y10VDD X115Y10VDD 25mOhm
L_X110Y10VDD_X120Y10VDD X115Y10VDD X120Y10VDD 2.91e-06nH
R_X110Y10VSS_X120Y10VSS X110Y10VSS X115Y10VSS 25mOhm
L_X110Y10VSS_X120Y10VSS X115Y10VSS X120Y10VSS 2.91e-06nH
R_X10Y20VDD_X20Y20VDD X10Y20VDD X15Y20VDD 25mOhm
L_X10Y20VDD_X20Y20VDD X15Y20VDD X20Y20VDD 2.91e-06nH
R_X10Y20VSS_X20Y20VSS X10Y20VSS X15Y20VSS 25mOhm
L_X10Y20VSS_X20Y20VSS X15Y20VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X30Y20VDD X20Y20VDD X25Y20VDD 25mOhm
L_X20Y20VDD_X30Y20VDD X25Y20VDD X30Y20VDD 2.91e-06nH
R_X20Y20VSS_X30Y20VSS X20Y20VSS X25Y20VSS 25mOhm
L_X20Y20VSS_X30Y20VSS X25Y20VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X40Y20VDD X30Y20VDD X35Y20VDD 25mOhm
L_X30Y20VDD_X40Y20VDD X35Y20VDD X40Y20VDD 2.91e-06nH
R_X30Y20VSS_X40Y20VSS X30Y20VSS X35Y20VSS 25mOhm
L_X30Y20VSS_X40Y20VSS X35Y20VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X50Y20VDD X40Y20VDD X45Y20VDD 25mOhm
L_X40Y20VDD_X50Y20VDD X45Y20VDD X50Y20VDD 2.91e-06nH
R_X40Y20VSS_X50Y20VSS X40Y20VSS X45Y20VSS 25mOhm
L_X40Y20VSS_X50Y20VSS X45Y20VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X60Y20VDD X50Y20VDD X55Y20VDD 25mOhm
L_X50Y20VDD_X60Y20VDD X55Y20VDD X60Y20VDD 2.91e-06nH
R_X50Y20VSS_X60Y20VSS X50Y20VSS X55Y20VSS 25mOhm
L_X50Y20VSS_X60Y20VSS X55Y20VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X70Y20VDD X60Y20VDD X65Y20VDD 25mOhm
L_X60Y20VDD_X70Y20VDD X65Y20VDD X70Y20VDD 2.91e-06nH
R_X60Y20VSS_X70Y20VSS X60Y20VSS X65Y20VSS 25mOhm
L_X60Y20VSS_X70Y20VSS X65Y20VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X80Y20VDD X70Y20VDD X75Y20VDD 25mOhm
L_X70Y20VDD_X80Y20VDD X75Y20VDD X80Y20VDD 2.91e-06nH
R_X70Y20VSS_X80Y20VSS X70Y20VSS X75Y20VSS 25mOhm
L_X70Y20VSS_X80Y20VSS X75Y20VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X90Y20VDD X80Y20VDD X85Y20VDD 25mOhm
L_X80Y20VDD_X90Y20VDD X85Y20VDD X90Y20VDD 2.91e-06nH
R_X80Y20VSS_X90Y20VSS X80Y20VSS X85Y20VSS 25mOhm
L_X80Y20VSS_X90Y20VSS X85Y20VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X100Y20VDD X90Y20VDD X95Y20VDD 25mOhm
L_X90Y20VDD_X100Y20VDD X95Y20VDD X100Y20VDD 2.91e-06nH
R_X90Y20VSS_X100Y20VSS X90Y20VSS X95Y20VSS 25mOhm
L_X90Y20VSS_X100Y20VSS X95Y20VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X110Y20VDD X100Y20VDD X105Y20VDD 25mOhm
L_X100Y20VDD_X110Y20VDD X105Y20VDD X110Y20VDD 2.91e-06nH
R_X100Y20VSS_X110Y20VSS X100Y20VSS X105Y20VSS 25mOhm
L_X100Y20VSS_X110Y20VSS X105Y20VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X120Y20VDD X110Y20VDD X115Y20VDD 25mOhm
L_X110Y20VDD_X120Y20VDD X115Y20VDD X120Y20VDD 2.91e-06nH
R_X110Y20VSS_X120Y20VSS X110Y20VSS X115Y20VSS 25mOhm
L_X110Y20VSS_X120Y20VSS X115Y20VSS X120Y20VSS 2.91e-06nH
R_X10Y30VDD_X20Y30VDD X10Y30VDD X15Y30VDD 25mOhm
L_X10Y30VDD_X20Y30VDD X15Y30VDD X20Y30VDD 2.91e-06nH
R_X10Y30VSS_X20Y30VSS X10Y30VSS X15Y30VSS 25mOhm
L_X10Y30VSS_X20Y30VSS X15Y30VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X30Y30VDD X20Y30VDD X25Y30VDD 25mOhm
L_X20Y30VDD_X30Y30VDD X25Y30VDD X30Y30VDD 2.91e-06nH
R_X20Y30VSS_X30Y30VSS X20Y30VSS X25Y30VSS 25mOhm
L_X20Y30VSS_X30Y30VSS X25Y30VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X40Y30VDD X30Y30VDD X35Y30VDD 25mOhm
L_X30Y30VDD_X40Y30VDD X35Y30VDD X40Y30VDD 2.91e-06nH
R_X30Y30VSS_X40Y30VSS X30Y30VSS X35Y30VSS 25mOhm
L_X30Y30VSS_X40Y30VSS X35Y30VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X50Y30VDD X40Y30VDD X45Y30VDD 25mOhm
L_X40Y30VDD_X50Y30VDD X45Y30VDD X50Y30VDD 2.91e-06nH
R_X40Y30VSS_X50Y30VSS X40Y30VSS X45Y30VSS 25mOhm
L_X40Y30VSS_X50Y30VSS X45Y30VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X60Y30VDD X50Y30VDD X55Y30VDD 25mOhm
L_X50Y30VDD_X60Y30VDD X55Y30VDD X60Y30VDD 2.91e-06nH
R_X50Y30VSS_X60Y30VSS X50Y30VSS X55Y30VSS 25mOhm
L_X50Y30VSS_X60Y30VSS X55Y30VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X70Y30VDD X60Y30VDD X65Y30VDD 25mOhm
L_X60Y30VDD_X70Y30VDD X65Y30VDD X70Y30VDD 2.91e-06nH
R_X60Y30VSS_X70Y30VSS X60Y30VSS X65Y30VSS 25mOhm
L_X60Y30VSS_X70Y30VSS X65Y30VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X80Y30VDD X70Y30VDD X75Y30VDD 25mOhm
L_X70Y30VDD_X80Y30VDD X75Y30VDD X80Y30VDD 2.91e-06nH
R_X70Y30VSS_X80Y30VSS X70Y30VSS X75Y30VSS 25mOhm
L_X70Y30VSS_X80Y30VSS X75Y30VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X90Y30VDD X80Y30VDD X85Y30VDD 25mOhm
L_X80Y30VDD_X90Y30VDD X85Y30VDD X90Y30VDD 2.91e-06nH
R_X80Y30VSS_X90Y30VSS X80Y30VSS X85Y30VSS 25mOhm
L_X80Y30VSS_X90Y30VSS X85Y30VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X100Y30VDD X90Y30VDD X95Y30VDD 25mOhm
L_X90Y30VDD_X100Y30VDD X95Y30VDD X100Y30VDD 2.91e-06nH
R_X90Y30VSS_X100Y30VSS X90Y30VSS X95Y30VSS 25mOhm
L_X90Y30VSS_X100Y30VSS X95Y30VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X110Y30VDD X100Y30VDD X105Y30VDD 25mOhm
L_X100Y30VDD_X110Y30VDD X105Y30VDD X110Y30VDD 2.91e-06nH
R_X100Y30VSS_X110Y30VSS X100Y30VSS X105Y30VSS 25mOhm
L_X100Y30VSS_X110Y30VSS X105Y30VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X120Y30VDD X110Y30VDD X115Y30VDD 25mOhm
L_X110Y30VDD_X120Y30VDD X115Y30VDD X120Y30VDD 2.91e-06nH
R_X110Y30VSS_X120Y30VSS X110Y30VSS X115Y30VSS 25mOhm
L_X110Y30VSS_X120Y30VSS X115Y30VSS X120Y30VSS 2.91e-06nH
R_X10Y40VDD_X20Y40VDD X10Y40VDD X15Y40VDD 25mOhm
L_X10Y40VDD_X20Y40VDD X15Y40VDD X20Y40VDD 2.91e-06nH
R_X10Y40VSS_X20Y40VSS X10Y40VSS X15Y40VSS 25mOhm
L_X10Y40VSS_X20Y40VSS X15Y40VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X30Y40VDD X20Y40VDD X25Y40VDD 25mOhm
L_X20Y40VDD_X30Y40VDD X25Y40VDD X30Y40VDD 2.91e-06nH
R_X20Y40VSS_X30Y40VSS X20Y40VSS X25Y40VSS 25mOhm
L_X20Y40VSS_X30Y40VSS X25Y40VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X40Y40VDD X30Y40VDD X35Y40VDD 25mOhm
L_X30Y40VDD_X40Y40VDD X35Y40VDD X40Y40VDD 2.91e-06nH
R_X30Y40VSS_X40Y40VSS X30Y40VSS X35Y40VSS 25mOhm
L_X30Y40VSS_X40Y40VSS X35Y40VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X50Y40VDD X40Y40VDD X45Y40VDD 25mOhm
L_X40Y40VDD_X50Y40VDD X45Y40VDD X50Y40VDD 2.91e-06nH
R_X40Y40VSS_X50Y40VSS X40Y40VSS X45Y40VSS 25mOhm
L_X40Y40VSS_X50Y40VSS X45Y40VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X60Y40VDD X50Y40VDD X55Y40VDD 25mOhm
L_X50Y40VDD_X60Y40VDD X55Y40VDD X60Y40VDD 2.91e-06nH
R_X50Y40VSS_X60Y40VSS X50Y40VSS X55Y40VSS 25mOhm
L_X50Y40VSS_X60Y40VSS X55Y40VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X70Y40VDD X60Y40VDD X65Y40VDD 25mOhm
L_X60Y40VDD_X70Y40VDD X65Y40VDD X70Y40VDD 2.91e-06nH
R_X60Y40VSS_X70Y40VSS X60Y40VSS X65Y40VSS 25mOhm
L_X60Y40VSS_X70Y40VSS X65Y40VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X80Y40VDD X70Y40VDD X75Y40VDD 25mOhm
L_X70Y40VDD_X80Y40VDD X75Y40VDD X80Y40VDD 2.91e-06nH
R_X70Y40VSS_X80Y40VSS X70Y40VSS X75Y40VSS 25mOhm
L_X70Y40VSS_X80Y40VSS X75Y40VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X90Y40VDD X80Y40VDD X85Y40VDD 25mOhm
L_X80Y40VDD_X90Y40VDD X85Y40VDD X90Y40VDD 2.91e-06nH
R_X80Y40VSS_X90Y40VSS X80Y40VSS X85Y40VSS 25mOhm
L_X80Y40VSS_X90Y40VSS X85Y40VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X100Y40VDD X90Y40VDD X95Y40VDD 25mOhm
L_X90Y40VDD_X100Y40VDD X95Y40VDD X100Y40VDD 2.91e-06nH
R_X90Y40VSS_X100Y40VSS X90Y40VSS X95Y40VSS 25mOhm
L_X90Y40VSS_X100Y40VSS X95Y40VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X110Y40VDD X100Y40VDD X105Y40VDD 25mOhm
L_X100Y40VDD_X110Y40VDD X105Y40VDD X110Y40VDD 2.91e-06nH
R_X100Y40VSS_X110Y40VSS X100Y40VSS X105Y40VSS 25mOhm
L_X100Y40VSS_X110Y40VSS X105Y40VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X120Y40VDD X110Y40VDD X115Y40VDD 25mOhm
L_X110Y40VDD_X120Y40VDD X115Y40VDD X120Y40VDD 2.91e-06nH
R_X110Y40VSS_X120Y40VSS X110Y40VSS X115Y40VSS 25mOhm
L_X110Y40VSS_X120Y40VSS X115Y40VSS X120Y40VSS 2.91e-06nH
R_X10Y50VDD_X20Y50VDD X10Y50VDD X15Y50VDD 25mOhm
L_X10Y50VDD_X20Y50VDD X15Y50VDD X20Y50VDD 2.91e-06nH
R_X10Y50VSS_X20Y50VSS X10Y50VSS X15Y50VSS 25mOhm
L_X10Y50VSS_X20Y50VSS X15Y50VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X30Y50VDD X20Y50VDD X25Y50VDD 25mOhm
L_X20Y50VDD_X30Y50VDD X25Y50VDD X30Y50VDD 2.91e-06nH
R_X20Y50VSS_X30Y50VSS X20Y50VSS X25Y50VSS 25mOhm
L_X20Y50VSS_X30Y50VSS X25Y50VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X40Y50VDD X30Y50VDD X35Y50VDD 25mOhm
L_X30Y50VDD_X40Y50VDD X35Y50VDD X40Y50VDD 2.91e-06nH
R_X30Y50VSS_X40Y50VSS X30Y50VSS X35Y50VSS 25mOhm
L_X30Y50VSS_X40Y50VSS X35Y50VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X50Y50VDD X40Y50VDD X45Y50VDD 25mOhm
L_X40Y50VDD_X50Y50VDD X45Y50VDD X50Y50VDD 2.91e-06nH
R_X40Y50VSS_X50Y50VSS X40Y50VSS X45Y50VSS 25mOhm
L_X40Y50VSS_X50Y50VSS X45Y50VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X60Y50VDD X50Y50VDD X55Y50VDD 25mOhm
L_X50Y50VDD_X60Y50VDD X55Y50VDD X60Y50VDD 2.91e-06nH
R_X50Y50VSS_X60Y50VSS X50Y50VSS X55Y50VSS 25mOhm
L_X50Y50VSS_X60Y50VSS X55Y50VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X70Y50VDD X60Y50VDD X65Y50VDD 25mOhm
L_X60Y50VDD_X70Y50VDD X65Y50VDD X70Y50VDD 2.91e-06nH
R_X60Y50VSS_X70Y50VSS X60Y50VSS X65Y50VSS 25mOhm
L_X60Y50VSS_X70Y50VSS X65Y50VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X80Y50VDD X70Y50VDD X75Y50VDD 25mOhm
L_X70Y50VDD_X80Y50VDD X75Y50VDD X80Y50VDD 2.91e-06nH
R_X70Y50VSS_X80Y50VSS X70Y50VSS X75Y50VSS 25mOhm
L_X70Y50VSS_X80Y50VSS X75Y50VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X90Y50VDD X80Y50VDD X85Y50VDD 25mOhm
L_X80Y50VDD_X90Y50VDD X85Y50VDD X90Y50VDD 2.91e-06nH
R_X80Y50VSS_X90Y50VSS X80Y50VSS X85Y50VSS 25mOhm
L_X80Y50VSS_X90Y50VSS X85Y50VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X100Y50VDD X90Y50VDD X95Y50VDD 25mOhm
L_X90Y50VDD_X100Y50VDD X95Y50VDD X100Y50VDD 2.91e-06nH
R_X90Y50VSS_X100Y50VSS X90Y50VSS X95Y50VSS 25mOhm
L_X90Y50VSS_X100Y50VSS X95Y50VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X110Y50VDD X100Y50VDD X105Y50VDD 25mOhm
L_X100Y50VDD_X110Y50VDD X105Y50VDD X110Y50VDD 2.91e-06nH
R_X100Y50VSS_X110Y50VSS X100Y50VSS X105Y50VSS 25mOhm
L_X100Y50VSS_X110Y50VSS X105Y50VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X120Y50VDD X110Y50VDD X115Y50VDD 25mOhm
L_X110Y50VDD_X120Y50VDD X115Y50VDD X120Y50VDD 2.91e-06nH
R_X110Y50VSS_X120Y50VSS X110Y50VSS X115Y50VSS 25mOhm
L_X110Y50VSS_X120Y50VSS X115Y50VSS X120Y50VSS 2.91e-06nH
R_X10Y60VDD_X20Y60VDD X10Y60VDD X15Y60VDD 25mOhm
L_X10Y60VDD_X20Y60VDD X15Y60VDD X20Y60VDD 2.91e-06nH
R_X10Y60VSS_X20Y60VSS X10Y60VSS X15Y60VSS 25mOhm
L_X10Y60VSS_X20Y60VSS X15Y60VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X30Y60VDD X20Y60VDD X25Y60VDD 25mOhm
L_X20Y60VDD_X30Y60VDD X25Y60VDD X30Y60VDD 2.91e-06nH
R_X20Y60VSS_X30Y60VSS X20Y60VSS X25Y60VSS 25mOhm
L_X20Y60VSS_X30Y60VSS X25Y60VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X40Y60VDD X30Y60VDD X35Y60VDD 25mOhm
L_X30Y60VDD_X40Y60VDD X35Y60VDD X40Y60VDD 2.91e-06nH
R_X30Y60VSS_X40Y60VSS X30Y60VSS X35Y60VSS 25mOhm
L_X30Y60VSS_X40Y60VSS X35Y60VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X50Y60VDD X40Y60VDD X45Y60VDD 25mOhm
L_X40Y60VDD_X50Y60VDD X45Y60VDD X50Y60VDD 2.91e-06nH
R_X40Y60VSS_X50Y60VSS X40Y60VSS X45Y60VSS 25mOhm
L_X40Y60VSS_X50Y60VSS X45Y60VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X60Y60VDD X50Y60VDD X55Y60VDD 25mOhm
L_X50Y60VDD_X60Y60VDD X55Y60VDD X60Y60VDD 2.91e-06nH
R_X50Y60VSS_X60Y60VSS X50Y60VSS X55Y60VSS 25mOhm
L_X50Y60VSS_X60Y60VSS X55Y60VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X70Y60VDD X60Y60VDD X65Y60VDD 25mOhm
L_X60Y60VDD_X70Y60VDD X65Y60VDD X70Y60VDD 2.91e-06nH
R_X60Y60VSS_X70Y60VSS X60Y60VSS X65Y60VSS 25mOhm
L_X60Y60VSS_X70Y60VSS X65Y60VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X80Y60VDD X70Y60VDD X75Y60VDD 25mOhm
L_X70Y60VDD_X80Y60VDD X75Y60VDD X80Y60VDD 2.91e-06nH
R_X70Y60VSS_X80Y60VSS X70Y60VSS X75Y60VSS 25mOhm
L_X70Y60VSS_X80Y60VSS X75Y60VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X90Y60VDD X80Y60VDD X85Y60VDD 25mOhm
L_X80Y60VDD_X90Y60VDD X85Y60VDD X90Y60VDD 2.91e-06nH
R_X80Y60VSS_X90Y60VSS X80Y60VSS X85Y60VSS 25mOhm
L_X80Y60VSS_X90Y60VSS X85Y60VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X100Y60VDD X90Y60VDD X95Y60VDD 25mOhm
L_X90Y60VDD_X100Y60VDD X95Y60VDD X100Y60VDD 2.91e-06nH
R_X90Y60VSS_X100Y60VSS X90Y60VSS X95Y60VSS 25mOhm
L_X90Y60VSS_X100Y60VSS X95Y60VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X110Y60VDD X100Y60VDD X105Y60VDD 25mOhm
L_X100Y60VDD_X110Y60VDD X105Y60VDD X110Y60VDD 2.91e-06nH
R_X100Y60VSS_X110Y60VSS X100Y60VSS X105Y60VSS 25mOhm
L_X100Y60VSS_X110Y60VSS X105Y60VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X120Y60VDD X110Y60VDD X115Y60VDD 25mOhm
L_X110Y60VDD_X120Y60VDD X115Y60VDD X120Y60VDD 2.91e-06nH
R_X110Y60VSS_X120Y60VSS X110Y60VSS X115Y60VSS 25mOhm
L_X110Y60VSS_X120Y60VSS X115Y60VSS X120Y60VSS 2.91e-06nH
R_X10Y70VDD_X20Y70VDD X10Y70VDD X15Y70VDD 25mOhm
L_X10Y70VDD_X20Y70VDD X15Y70VDD X20Y70VDD 2.91e-06nH
R_X10Y70VSS_X20Y70VSS X10Y70VSS X15Y70VSS 25mOhm
L_X10Y70VSS_X20Y70VSS X15Y70VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X30Y70VDD X20Y70VDD X25Y70VDD 25mOhm
L_X20Y70VDD_X30Y70VDD X25Y70VDD X30Y70VDD 2.91e-06nH
R_X20Y70VSS_X30Y70VSS X20Y70VSS X25Y70VSS 25mOhm
L_X20Y70VSS_X30Y70VSS X25Y70VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X40Y70VDD X30Y70VDD X35Y70VDD 25mOhm
L_X30Y70VDD_X40Y70VDD X35Y70VDD X40Y70VDD 2.91e-06nH
R_X30Y70VSS_X40Y70VSS X30Y70VSS X35Y70VSS 25mOhm
L_X30Y70VSS_X40Y70VSS X35Y70VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X50Y70VDD X40Y70VDD X45Y70VDD 25mOhm
L_X40Y70VDD_X50Y70VDD X45Y70VDD X50Y70VDD 2.91e-06nH
R_X40Y70VSS_X50Y70VSS X40Y70VSS X45Y70VSS 25mOhm
L_X40Y70VSS_X50Y70VSS X45Y70VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X60Y70VDD X50Y70VDD X55Y70VDD 25mOhm
L_X50Y70VDD_X60Y70VDD X55Y70VDD X60Y70VDD 2.91e-06nH
R_X50Y70VSS_X60Y70VSS X50Y70VSS X55Y70VSS 25mOhm
L_X50Y70VSS_X60Y70VSS X55Y70VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X70Y70VDD X60Y70VDD X65Y70VDD 25mOhm
L_X60Y70VDD_X70Y70VDD X65Y70VDD X70Y70VDD 2.91e-06nH
R_X60Y70VSS_X70Y70VSS X60Y70VSS X65Y70VSS 25mOhm
L_X60Y70VSS_X70Y70VSS X65Y70VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X80Y70VDD X70Y70VDD X75Y70VDD 25mOhm
L_X70Y70VDD_X80Y70VDD X75Y70VDD X80Y70VDD 2.91e-06nH
R_X70Y70VSS_X80Y70VSS X70Y70VSS X75Y70VSS 25mOhm
L_X70Y70VSS_X80Y70VSS X75Y70VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X90Y70VDD X80Y70VDD X85Y70VDD 25mOhm
L_X80Y70VDD_X90Y70VDD X85Y70VDD X90Y70VDD 2.91e-06nH
R_X80Y70VSS_X90Y70VSS X80Y70VSS X85Y70VSS 25mOhm
L_X80Y70VSS_X90Y70VSS X85Y70VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X100Y70VDD X90Y70VDD X95Y70VDD 25mOhm
L_X90Y70VDD_X100Y70VDD X95Y70VDD X100Y70VDD 2.91e-06nH
R_X90Y70VSS_X100Y70VSS X90Y70VSS X95Y70VSS 25mOhm
L_X90Y70VSS_X100Y70VSS X95Y70VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X110Y70VDD X100Y70VDD X105Y70VDD 25mOhm
L_X100Y70VDD_X110Y70VDD X105Y70VDD X110Y70VDD 2.91e-06nH
R_X100Y70VSS_X110Y70VSS X100Y70VSS X105Y70VSS 25mOhm
L_X100Y70VSS_X110Y70VSS X105Y70VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X120Y70VDD X110Y70VDD X115Y70VDD 25mOhm
L_X110Y70VDD_X120Y70VDD X115Y70VDD X120Y70VDD 2.91e-06nH
R_X110Y70VSS_X120Y70VSS X110Y70VSS X115Y70VSS 25mOhm
L_X110Y70VSS_X120Y70VSS X115Y70VSS X120Y70VSS 2.91e-06nH
R_X10Y80VDD_X20Y80VDD X10Y80VDD X15Y80VDD 25mOhm
L_X10Y80VDD_X20Y80VDD X15Y80VDD X20Y80VDD 2.91e-06nH
R_X10Y80VSS_X20Y80VSS X10Y80VSS X15Y80VSS 25mOhm
L_X10Y80VSS_X20Y80VSS X15Y80VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X30Y80VDD X20Y80VDD X25Y80VDD 25mOhm
L_X20Y80VDD_X30Y80VDD X25Y80VDD X30Y80VDD 2.91e-06nH
R_X20Y80VSS_X30Y80VSS X20Y80VSS X25Y80VSS 25mOhm
L_X20Y80VSS_X30Y80VSS X25Y80VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X40Y80VDD X30Y80VDD X35Y80VDD 25mOhm
L_X30Y80VDD_X40Y80VDD X35Y80VDD X40Y80VDD 2.91e-06nH
R_X30Y80VSS_X40Y80VSS X30Y80VSS X35Y80VSS 25mOhm
L_X30Y80VSS_X40Y80VSS X35Y80VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X50Y80VDD X40Y80VDD X45Y80VDD 25mOhm
L_X40Y80VDD_X50Y80VDD X45Y80VDD X50Y80VDD 2.91e-06nH
R_X40Y80VSS_X50Y80VSS X40Y80VSS X45Y80VSS 25mOhm
L_X40Y80VSS_X50Y80VSS X45Y80VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X60Y80VDD X50Y80VDD X55Y80VDD 25mOhm
L_X50Y80VDD_X60Y80VDD X55Y80VDD X60Y80VDD 2.91e-06nH
R_X50Y80VSS_X60Y80VSS X50Y80VSS X55Y80VSS 25mOhm
L_X50Y80VSS_X60Y80VSS X55Y80VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X70Y80VDD X60Y80VDD X65Y80VDD 25mOhm
L_X60Y80VDD_X70Y80VDD X65Y80VDD X70Y80VDD 2.91e-06nH
R_X60Y80VSS_X70Y80VSS X60Y80VSS X65Y80VSS 25mOhm
L_X60Y80VSS_X70Y80VSS X65Y80VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X80Y80VDD X70Y80VDD X75Y80VDD 25mOhm
L_X70Y80VDD_X80Y80VDD X75Y80VDD X80Y80VDD 2.91e-06nH
R_X70Y80VSS_X80Y80VSS X70Y80VSS X75Y80VSS 25mOhm
L_X70Y80VSS_X80Y80VSS X75Y80VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X90Y80VDD X80Y80VDD X85Y80VDD 25mOhm
L_X80Y80VDD_X90Y80VDD X85Y80VDD X90Y80VDD 2.91e-06nH
R_X80Y80VSS_X90Y80VSS X80Y80VSS X85Y80VSS 25mOhm
L_X80Y80VSS_X90Y80VSS X85Y80VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X100Y80VDD X90Y80VDD X95Y80VDD 25mOhm
L_X90Y80VDD_X100Y80VDD X95Y80VDD X100Y80VDD 2.91e-06nH
R_X90Y80VSS_X100Y80VSS X90Y80VSS X95Y80VSS 25mOhm
L_X90Y80VSS_X100Y80VSS X95Y80VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X110Y80VDD X100Y80VDD X105Y80VDD 25mOhm
L_X100Y80VDD_X110Y80VDD X105Y80VDD X110Y80VDD 2.91e-06nH
R_X100Y80VSS_X110Y80VSS X100Y80VSS X105Y80VSS 25mOhm
L_X100Y80VSS_X110Y80VSS X105Y80VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X120Y80VDD X110Y80VDD X115Y80VDD 25mOhm
L_X110Y80VDD_X120Y80VDD X115Y80VDD X120Y80VDD 2.91e-06nH
R_X110Y80VSS_X120Y80VSS X110Y80VSS X115Y80VSS 25mOhm
L_X110Y80VSS_X120Y80VSS X115Y80VSS X120Y80VSS 2.91e-06nH
R_X10Y90VDD_X20Y90VDD X10Y90VDD X15Y90VDD 25mOhm
L_X10Y90VDD_X20Y90VDD X15Y90VDD X20Y90VDD 2.91e-06nH
R_X10Y90VSS_X20Y90VSS X10Y90VSS X15Y90VSS 25mOhm
L_X10Y90VSS_X20Y90VSS X15Y90VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X30Y90VDD X20Y90VDD X25Y90VDD 25mOhm
L_X20Y90VDD_X30Y90VDD X25Y90VDD X30Y90VDD 2.91e-06nH
R_X20Y90VSS_X30Y90VSS X20Y90VSS X25Y90VSS 25mOhm
L_X20Y90VSS_X30Y90VSS X25Y90VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X40Y90VDD X30Y90VDD X35Y90VDD 25mOhm
L_X30Y90VDD_X40Y90VDD X35Y90VDD X40Y90VDD 2.91e-06nH
R_X30Y90VSS_X40Y90VSS X30Y90VSS X35Y90VSS 25mOhm
L_X30Y90VSS_X40Y90VSS X35Y90VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X50Y90VDD X40Y90VDD X45Y90VDD 25mOhm
L_X40Y90VDD_X50Y90VDD X45Y90VDD X50Y90VDD 2.91e-06nH
R_X40Y90VSS_X50Y90VSS X40Y90VSS X45Y90VSS 25mOhm
L_X40Y90VSS_X50Y90VSS X45Y90VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X60Y90VDD X50Y90VDD X55Y90VDD 25mOhm
L_X50Y90VDD_X60Y90VDD X55Y90VDD X60Y90VDD 2.91e-06nH
R_X50Y90VSS_X60Y90VSS X50Y90VSS X55Y90VSS 25mOhm
L_X50Y90VSS_X60Y90VSS X55Y90VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X70Y90VDD X60Y90VDD X65Y90VDD 25mOhm
L_X60Y90VDD_X70Y90VDD X65Y90VDD X70Y90VDD 2.91e-06nH
R_X60Y90VSS_X70Y90VSS X60Y90VSS X65Y90VSS 25mOhm
L_X60Y90VSS_X70Y90VSS X65Y90VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X80Y90VDD X70Y90VDD X75Y90VDD 25mOhm
L_X70Y90VDD_X80Y90VDD X75Y90VDD X80Y90VDD 2.91e-06nH
R_X70Y90VSS_X80Y90VSS X70Y90VSS X75Y90VSS 25mOhm
L_X70Y90VSS_X80Y90VSS X75Y90VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X90Y90VDD X80Y90VDD X85Y90VDD 25mOhm
L_X80Y90VDD_X90Y90VDD X85Y90VDD X90Y90VDD 2.91e-06nH
R_X80Y90VSS_X90Y90VSS X80Y90VSS X85Y90VSS 25mOhm
L_X80Y90VSS_X90Y90VSS X85Y90VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X100Y90VDD X90Y90VDD X95Y90VDD 25mOhm
L_X90Y90VDD_X100Y90VDD X95Y90VDD X100Y90VDD 2.91e-06nH
R_X90Y90VSS_X100Y90VSS X90Y90VSS X95Y90VSS 25mOhm
L_X90Y90VSS_X100Y90VSS X95Y90VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X110Y90VDD X100Y90VDD X105Y90VDD 25mOhm
L_X100Y90VDD_X110Y90VDD X105Y90VDD X110Y90VDD 2.91e-06nH
R_X100Y90VSS_X110Y90VSS X100Y90VSS X105Y90VSS 25mOhm
L_X100Y90VSS_X110Y90VSS X105Y90VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X120Y90VDD X110Y90VDD X115Y90VDD 25mOhm
L_X110Y90VDD_X120Y90VDD X115Y90VDD X120Y90VDD 2.91e-06nH
R_X110Y90VSS_X120Y90VSS X110Y90VSS X115Y90VSS 25mOhm
L_X110Y90VSS_X120Y90VSS X115Y90VSS X120Y90VSS 2.91e-06nH
R_X10Y100VDD_X20Y100VDD X10Y100VDD X15Y100VDD 25mOhm
L_X10Y100VDD_X20Y100VDD X15Y100VDD X20Y100VDD 2.91e-06nH
R_X10Y100VSS_X20Y100VSS X10Y100VSS X15Y100VSS 25mOhm
L_X10Y100VSS_X20Y100VSS X15Y100VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X30Y100VDD X20Y100VDD X25Y100VDD 25mOhm
L_X20Y100VDD_X30Y100VDD X25Y100VDD X30Y100VDD 2.91e-06nH
R_X20Y100VSS_X30Y100VSS X20Y100VSS X25Y100VSS 25mOhm
L_X20Y100VSS_X30Y100VSS X25Y100VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X40Y100VDD X30Y100VDD X35Y100VDD 25mOhm
L_X30Y100VDD_X40Y100VDD X35Y100VDD X40Y100VDD 2.91e-06nH
R_X30Y100VSS_X40Y100VSS X30Y100VSS X35Y100VSS 25mOhm
L_X30Y100VSS_X40Y100VSS X35Y100VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X50Y100VDD X40Y100VDD X45Y100VDD 25mOhm
L_X40Y100VDD_X50Y100VDD X45Y100VDD X50Y100VDD 2.91e-06nH
R_X40Y100VSS_X50Y100VSS X40Y100VSS X45Y100VSS 25mOhm
L_X40Y100VSS_X50Y100VSS X45Y100VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X60Y100VDD X50Y100VDD X55Y100VDD 25mOhm
L_X50Y100VDD_X60Y100VDD X55Y100VDD X60Y100VDD 2.91e-06nH
R_X50Y100VSS_X60Y100VSS X50Y100VSS X55Y100VSS 25mOhm
L_X50Y100VSS_X60Y100VSS X55Y100VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X70Y100VDD X60Y100VDD X65Y100VDD 25mOhm
L_X60Y100VDD_X70Y100VDD X65Y100VDD X70Y100VDD 2.91e-06nH
R_X60Y100VSS_X70Y100VSS X60Y100VSS X65Y100VSS 25mOhm
L_X60Y100VSS_X70Y100VSS X65Y100VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X80Y100VDD X70Y100VDD X75Y100VDD 25mOhm
L_X70Y100VDD_X80Y100VDD X75Y100VDD X80Y100VDD 2.91e-06nH
R_X70Y100VSS_X80Y100VSS X70Y100VSS X75Y100VSS 25mOhm
L_X70Y100VSS_X80Y100VSS X75Y100VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X90Y100VDD X80Y100VDD X85Y100VDD 25mOhm
L_X80Y100VDD_X90Y100VDD X85Y100VDD X90Y100VDD 2.91e-06nH
R_X80Y100VSS_X90Y100VSS X80Y100VSS X85Y100VSS 25mOhm
L_X80Y100VSS_X90Y100VSS X85Y100VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X100Y100VDD X90Y100VDD X95Y100VDD 25mOhm
L_X90Y100VDD_X100Y100VDD X95Y100VDD X100Y100VDD 2.91e-06nH
R_X90Y100VSS_X100Y100VSS X90Y100VSS X95Y100VSS 25mOhm
L_X90Y100VSS_X100Y100VSS X95Y100VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X110Y100VDD X100Y100VDD X105Y100VDD 25mOhm
L_X100Y100VDD_X110Y100VDD X105Y100VDD X110Y100VDD 2.91e-06nH
R_X100Y100VSS_X110Y100VSS X100Y100VSS X105Y100VSS 25mOhm
L_X100Y100VSS_X110Y100VSS X105Y100VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X120Y100VDD X110Y100VDD X115Y100VDD 25mOhm
L_X110Y100VDD_X120Y100VDD X115Y100VDD X120Y100VDD 2.91e-06nH
R_X110Y100VSS_X120Y100VSS X110Y100VSS X115Y100VSS 25mOhm
L_X110Y100VSS_X120Y100VSS X115Y100VSS X120Y100VSS 2.91e-06nH
R_X10Y110VDD_X20Y110VDD X10Y110VDD X15Y110VDD 25mOhm
L_X10Y110VDD_X20Y110VDD X15Y110VDD X20Y110VDD 2.91e-06nH
R_X10Y110VSS_X20Y110VSS X10Y110VSS X15Y110VSS 25mOhm
L_X10Y110VSS_X20Y110VSS X15Y110VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X30Y110VDD X20Y110VDD X25Y110VDD 25mOhm
L_X20Y110VDD_X30Y110VDD X25Y110VDD X30Y110VDD 2.91e-06nH
R_X20Y110VSS_X30Y110VSS X20Y110VSS X25Y110VSS 25mOhm
L_X20Y110VSS_X30Y110VSS X25Y110VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X40Y110VDD X30Y110VDD X35Y110VDD 25mOhm
L_X30Y110VDD_X40Y110VDD X35Y110VDD X40Y110VDD 2.91e-06nH
R_X30Y110VSS_X40Y110VSS X30Y110VSS X35Y110VSS 25mOhm
L_X30Y110VSS_X40Y110VSS X35Y110VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X50Y110VDD X40Y110VDD X45Y110VDD 25mOhm
L_X40Y110VDD_X50Y110VDD X45Y110VDD X50Y110VDD 2.91e-06nH
R_X40Y110VSS_X50Y110VSS X40Y110VSS X45Y110VSS 25mOhm
L_X40Y110VSS_X50Y110VSS X45Y110VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X60Y110VDD X50Y110VDD X55Y110VDD 25mOhm
L_X50Y110VDD_X60Y110VDD X55Y110VDD X60Y110VDD 2.91e-06nH
R_X50Y110VSS_X60Y110VSS X50Y110VSS X55Y110VSS 25mOhm
L_X50Y110VSS_X60Y110VSS X55Y110VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X70Y110VDD X60Y110VDD X65Y110VDD 25mOhm
L_X60Y110VDD_X70Y110VDD X65Y110VDD X70Y110VDD 2.91e-06nH
R_X60Y110VSS_X70Y110VSS X60Y110VSS X65Y110VSS 25mOhm
L_X60Y110VSS_X70Y110VSS X65Y110VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X80Y110VDD X70Y110VDD X75Y110VDD 25mOhm
L_X70Y110VDD_X80Y110VDD X75Y110VDD X80Y110VDD 2.91e-06nH
R_X70Y110VSS_X80Y110VSS X70Y110VSS X75Y110VSS 25mOhm
L_X70Y110VSS_X80Y110VSS X75Y110VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X90Y110VDD X80Y110VDD X85Y110VDD 25mOhm
L_X80Y110VDD_X90Y110VDD X85Y110VDD X90Y110VDD 2.91e-06nH
R_X80Y110VSS_X90Y110VSS X80Y110VSS X85Y110VSS 25mOhm
L_X80Y110VSS_X90Y110VSS X85Y110VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X100Y110VDD X90Y110VDD X95Y110VDD 25mOhm
L_X90Y110VDD_X100Y110VDD X95Y110VDD X100Y110VDD 2.91e-06nH
R_X90Y110VSS_X100Y110VSS X90Y110VSS X95Y110VSS 25mOhm
L_X90Y110VSS_X100Y110VSS X95Y110VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X110Y110VDD X100Y110VDD X105Y110VDD 25mOhm
L_X100Y110VDD_X110Y110VDD X105Y110VDD X110Y110VDD 2.91e-06nH
R_X100Y110VSS_X110Y110VSS X100Y110VSS X105Y110VSS 25mOhm
L_X100Y110VSS_X110Y110VSS X105Y110VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X120Y110VDD X110Y110VDD X115Y110VDD 25mOhm
L_X110Y110VDD_X120Y110VDD X115Y110VDD X120Y110VDD 2.91e-06nH
R_X110Y110VSS_X120Y110VSS X110Y110VSS X115Y110VSS 25mOhm
L_X110Y110VSS_X120Y110VSS X115Y110VSS X120Y110VSS 2.91e-06nH
R_X10Y120VDD_X20Y120VDD X10Y120VDD X15Y120VDD 25mOhm
L_X10Y120VDD_X20Y120VDD X15Y120VDD X20Y120VDD 2.91e-06nH
R_X10Y120VSS_X20Y120VSS X10Y120VSS X15Y120VSS 25mOhm
L_X10Y120VSS_X20Y120VSS X15Y120VSS X20Y120VSS 2.91e-06nH
R_X20Y120VDD_X30Y120VDD X20Y120VDD X25Y120VDD 25mOhm
L_X20Y120VDD_X30Y120VDD X25Y120VDD X30Y120VDD 2.91e-06nH
R_X20Y120VSS_X30Y120VSS X20Y120VSS X25Y120VSS 25mOhm
L_X20Y120VSS_X30Y120VSS X25Y120VSS X30Y120VSS 2.91e-06nH
R_X30Y120VDD_X40Y120VDD X30Y120VDD X35Y120VDD 25mOhm
L_X30Y120VDD_X40Y120VDD X35Y120VDD X40Y120VDD 2.91e-06nH
R_X30Y120VSS_X40Y120VSS X30Y120VSS X35Y120VSS 25mOhm
L_X30Y120VSS_X40Y120VSS X35Y120VSS X40Y120VSS 2.91e-06nH
R_X40Y120VDD_X50Y120VDD X40Y120VDD X45Y120VDD 25mOhm
L_X40Y120VDD_X50Y120VDD X45Y120VDD X50Y120VDD 2.91e-06nH
R_X40Y120VSS_X50Y120VSS X40Y120VSS X45Y120VSS 25mOhm
L_X40Y120VSS_X50Y120VSS X45Y120VSS X50Y120VSS 2.91e-06nH
R_X50Y120VDD_X60Y120VDD X50Y120VDD X55Y120VDD 25mOhm
L_X50Y120VDD_X60Y120VDD X55Y120VDD X60Y120VDD 2.91e-06nH
R_X50Y120VSS_X60Y120VSS X50Y120VSS X55Y120VSS 25mOhm
L_X50Y120VSS_X60Y120VSS X55Y120VSS X60Y120VSS 2.91e-06nH
R_X60Y120VDD_X70Y120VDD X60Y120VDD X65Y120VDD 25mOhm
L_X60Y120VDD_X70Y120VDD X65Y120VDD X70Y120VDD 2.91e-06nH
R_X60Y120VSS_X70Y120VSS X60Y120VSS X65Y120VSS 25mOhm
L_X60Y120VSS_X70Y120VSS X65Y120VSS X70Y120VSS 2.91e-06nH
R_X70Y120VDD_X80Y120VDD X70Y120VDD X75Y120VDD 25mOhm
L_X70Y120VDD_X80Y120VDD X75Y120VDD X80Y120VDD 2.91e-06nH
R_X70Y120VSS_X80Y120VSS X70Y120VSS X75Y120VSS 25mOhm
L_X70Y120VSS_X80Y120VSS X75Y120VSS X80Y120VSS 2.91e-06nH
R_X80Y120VDD_X90Y120VDD X80Y120VDD X85Y120VDD 25mOhm
L_X80Y120VDD_X90Y120VDD X85Y120VDD X90Y120VDD 2.91e-06nH
R_X80Y120VSS_X90Y120VSS X80Y120VSS X85Y120VSS 25mOhm
L_X80Y120VSS_X90Y120VSS X85Y120VSS X90Y120VSS 2.91e-06nH
R_X90Y120VDD_X100Y120VDD X90Y120VDD X95Y120VDD 25mOhm
L_X90Y120VDD_X100Y120VDD X95Y120VDD X100Y120VDD 2.91e-06nH
R_X90Y120VSS_X100Y120VSS X90Y120VSS X95Y120VSS 25mOhm
L_X90Y120VSS_X100Y120VSS X95Y120VSS X100Y120VSS 2.91e-06nH
R_X100Y120VDD_X110Y120VDD X100Y120VDD X105Y120VDD 25mOhm
L_X100Y120VDD_X110Y120VDD X105Y120VDD X110Y120VDD 2.91e-06nH
R_X100Y120VSS_X110Y120VSS X100Y120VSS X105Y120VSS 25mOhm
L_X100Y120VSS_X110Y120VSS X105Y120VSS X110Y120VSS 2.91e-06nH
R_X110Y120VDD_X120Y120VDD X110Y120VDD X115Y120VDD 25mOhm
L_X110Y120VDD_X120Y120VDD X115Y120VDD X120Y120VDD 2.91e-06nH
R_X110Y120VSS_X120Y120VSS X110Y120VSS X115Y120VSS 25mOhm
L_X110Y120VSS_X120Y120VSS X115Y120VSS X120Y120VSS 2.91e-06nH
R_X10Y10VDD_X10Y20VDD X10Y10VDD X10Y15VDD 25mOhm
L_X10Y10VDD_X10Y20VDD X10Y15VDD X10Y20VDD 2.91e-06nH
R_X10Y10VSS_X10Y20VSS X10Y10VSS X10Y15VSS 25mOhm
L_X10Y10VSS_X10Y20VSS X10Y15VSS X10Y20VSS 2.91e-06nH
R_X10Y20VDD_X10Y30VDD X10Y20VDD X10Y25VDD 25mOhm
L_X10Y20VDD_X10Y30VDD X10Y25VDD X10Y30VDD 2.91e-06nH
R_X10Y20VSS_X10Y30VSS X10Y20VSS X10Y25VSS 25mOhm
L_X10Y20VSS_X10Y30VSS X10Y25VSS X10Y30VSS 2.91e-06nH
R_X10Y30VDD_X10Y40VDD X10Y30VDD X10Y35VDD 25mOhm
L_X10Y30VDD_X10Y40VDD X10Y35VDD X10Y40VDD 2.91e-06nH
R_X10Y30VSS_X10Y40VSS X10Y30VSS X10Y35VSS 25mOhm
L_X10Y30VSS_X10Y40VSS X10Y35VSS X10Y40VSS 2.91e-06nH
R_X10Y40VDD_X10Y50VDD X10Y40VDD X10Y45VDD 25mOhm
L_X10Y40VDD_X10Y50VDD X10Y45VDD X10Y50VDD 2.91e-06nH
R_X10Y40VSS_X10Y50VSS X10Y40VSS X10Y45VSS 25mOhm
L_X10Y40VSS_X10Y50VSS X10Y45VSS X10Y50VSS 2.91e-06nH
R_X10Y50VDD_X10Y60VDD X10Y50VDD X10Y55VDD 25mOhm
L_X10Y50VDD_X10Y60VDD X10Y55VDD X10Y60VDD 2.91e-06nH
R_X10Y50VSS_X10Y60VSS X10Y50VSS X10Y55VSS 25mOhm
L_X10Y50VSS_X10Y60VSS X10Y55VSS X10Y60VSS 2.91e-06nH
R_X10Y60VDD_X10Y70VDD X10Y60VDD X10Y65VDD 25mOhm
L_X10Y60VDD_X10Y70VDD X10Y65VDD X10Y70VDD 2.91e-06nH
R_X10Y60VSS_X10Y70VSS X10Y60VSS X10Y65VSS 25mOhm
L_X10Y60VSS_X10Y70VSS X10Y65VSS X10Y70VSS 2.91e-06nH
R_X10Y70VDD_X10Y80VDD X10Y70VDD X10Y75VDD 25mOhm
L_X10Y70VDD_X10Y80VDD X10Y75VDD X10Y80VDD 2.91e-06nH
R_X10Y70VSS_X10Y80VSS X10Y70VSS X10Y75VSS 25mOhm
L_X10Y70VSS_X10Y80VSS X10Y75VSS X10Y80VSS 2.91e-06nH
R_X10Y80VDD_X10Y90VDD X10Y80VDD X10Y85VDD 25mOhm
L_X10Y80VDD_X10Y90VDD X10Y85VDD X10Y90VDD 2.91e-06nH
R_X10Y80VSS_X10Y90VSS X10Y80VSS X10Y85VSS 25mOhm
L_X10Y80VSS_X10Y90VSS X10Y85VSS X10Y90VSS 2.91e-06nH
R_X10Y90VDD_X10Y100VDD X10Y90VDD X10Y95VDD 25mOhm
L_X10Y90VDD_X10Y100VDD X10Y95VDD X10Y100VDD 2.91e-06nH
R_X10Y90VSS_X10Y100VSS X10Y90VSS X10Y95VSS 25mOhm
L_X10Y90VSS_X10Y100VSS X10Y95VSS X10Y100VSS 2.91e-06nH
R_X10Y100VDD_X10Y110VDD X10Y100VDD X10Y105VDD 25mOhm
L_X10Y100VDD_X10Y110VDD X10Y105VDD X10Y110VDD 2.91e-06nH
R_X10Y100VSS_X10Y110VSS X10Y100VSS X10Y105VSS 25mOhm
L_X10Y100VSS_X10Y110VSS X10Y105VSS X10Y110VSS 2.91e-06nH
R_X10Y110VDD_X10Y120VDD X10Y110VDD X10Y115VDD 25mOhm
L_X10Y110VDD_X10Y120VDD X10Y115VDD X10Y120VDD 2.91e-06nH
R_X10Y110VSS_X10Y120VSS X10Y110VSS X10Y115VSS 25mOhm
L_X10Y110VSS_X10Y120VSS X10Y115VSS X10Y120VSS 2.91e-06nH
R_X20Y10VDD_X20Y20VDD X20Y10VDD X20Y15VDD 25mOhm
L_X20Y10VDD_X20Y20VDD X20Y15VDD X20Y20VDD 2.91e-06nH
R_X20Y10VSS_X20Y20VSS X20Y10VSS X20Y15VSS 25mOhm
L_X20Y10VSS_X20Y20VSS X20Y15VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X20Y30VDD X20Y20VDD X20Y25VDD 25mOhm
L_X20Y20VDD_X20Y30VDD X20Y25VDD X20Y30VDD 2.91e-06nH
R_X20Y20VSS_X20Y30VSS X20Y20VSS X20Y25VSS 25mOhm
L_X20Y20VSS_X20Y30VSS X20Y25VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X20Y40VDD X20Y30VDD X20Y35VDD 25mOhm
L_X20Y30VDD_X20Y40VDD X20Y35VDD X20Y40VDD 2.91e-06nH
R_X20Y30VSS_X20Y40VSS X20Y30VSS X20Y35VSS 25mOhm
L_X20Y30VSS_X20Y40VSS X20Y35VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X20Y50VDD X20Y40VDD X20Y45VDD 25mOhm
L_X20Y40VDD_X20Y50VDD X20Y45VDD X20Y50VDD 2.91e-06nH
R_X20Y40VSS_X20Y50VSS X20Y40VSS X20Y45VSS 25mOhm
L_X20Y40VSS_X20Y50VSS X20Y45VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X20Y60VDD X20Y50VDD X20Y55VDD 25mOhm
L_X20Y50VDD_X20Y60VDD X20Y55VDD X20Y60VDD 2.91e-06nH
R_X20Y50VSS_X20Y60VSS X20Y50VSS X20Y55VSS 25mOhm
L_X20Y50VSS_X20Y60VSS X20Y55VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X20Y70VDD X20Y60VDD X20Y65VDD 25mOhm
L_X20Y60VDD_X20Y70VDD X20Y65VDD X20Y70VDD 2.91e-06nH
R_X20Y60VSS_X20Y70VSS X20Y60VSS X20Y65VSS 25mOhm
L_X20Y60VSS_X20Y70VSS X20Y65VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X20Y80VDD X20Y70VDD X20Y75VDD 25mOhm
L_X20Y70VDD_X20Y80VDD X20Y75VDD X20Y80VDD 2.91e-06nH
R_X20Y70VSS_X20Y80VSS X20Y70VSS X20Y75VSS 25mOhm
L_X20Y70VSS_X20Y80VSS X20Y75VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X20Y90VDD X20Y80VDD X20Y85VDD 25mOhm
L_X20Y80VDD_X20Y90VDD X20Y85VDD X20Y90VDD 2.91e-06nH
R_X20Y80VSS_X20Y90VSS X20Y80VSS X20Y85VSS 25mOhm
L_X20Y80VSS_X20Y90VSS X20Y85VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X20Y100VDD X20Y90VDD X20Y95VDD 25mOhm
L_X20Y90VDD_X20Y100VDD X20Y95VDD X20Y100VDD 2.91e-06nH
R_X20Y90VSS_X20Y100VSS X20Y90VSS X20Y95VSS 25mOhm
L_X20Y90VSS_X20Y100VSS X20Y95VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X20Y110VDD X20Y100VDD X20Y105VDD 25mOhm
L_X20Y100VDD_X20Y110VDD X20Y105VDD X20Y110VDD 2.91e-06nH
R_X20Y100VSS_X20Y110VSS X20Y100VSS X20Y105VSS 25mOhm
L_X20Y100VSS_X20Y110VSS X20Y105VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X20Y120VDD X20Y110VDD X20Y115VDD 25mOhm
L_X20Y110VDD_X20Y120VDD X20Y115VDD X20Y120VDD 2.91e-06nH
R_X20Y110VSS_X20Y120VSS X20Y110VSS X20Y115VSS 25mOhm
L_X20Y110VSS_X20Y120VSS X20Y115VSS X20Y120VSS 2.91e-06nH
R_X30Y10VDD_X30Y20VDD X30Y10VDD X30Y15VDD 25mOhm
L_X30Y10VDD_X30Y20VDD X30Y15VDD X30Y20VDD 2.91e-06nH
R_X30Y10VSS_X30Y20VSS X30Y10VSS X30Y15VSS 25mOhm
L_X30Y10VSS_X30Y20VSS X30Y15VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X30Y30VDD X30Y20VDD X30Y25VDD 25mOhm
L_X30Y20VDD_X30Y30VDD X30Y25VDD X30Y30VDD 2.91e-06nH
R_X30Y20VSS_X30Y30VSS X30Y20VSS X30Y25VSS 25mOhm
L_X30Y20VSS_X30Y30VSS X30Y25VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X30Y40VDD X30Y30VDD X30Y35VDD 25mOhm
L_X30Y30VDD_X30Y40VDD X30Y35VDD X30Y40VDD 2.91e-06nH
R_X30Y30VSS_X30Y40VSS X30Y30VSS X30Y35VSS 25mOhm
L_X30Y30VSS_X30Y40VSS X30Y35VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X30Y50VDD X30Y40VDD X30Y45VDD 25mOhm
L_X30Y40VDD_X30Y50VDD X30Y45VDD X30Y50VDD 2.91e-06nH
R_X30Y40VSS_X30Y50VSS X30Y40VSS X30Y45VSS 25mOhm
L_X30Y40VSS_X30Y50VSS X30Y45VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X30Y60VDD X30Y50VDD X30Y55VDD 25mOhm
L_X30Y50VDD_X30Y60VDD X30Y55VDD X30Y60VDD 2.91e-06nH
R_X30Y50VSS_X30Y60VSS X30Y50VSS X30Y55VSS 25mOhm
L_X30Y50VSS_X30Y60VSS X30Y55VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X30Y70VDD X30Y60VDD X30Y65VDD 25mOhm
L_X30Y60VDD_X30Y70VDD X30Y65VDD X30Y70VDD 2.91e-06nH
R_X30Y60VSS_X30Y70VSS X30Y60VSS X30Y65VSS 25mOhm
L_X30Y60VSS_X30Y70VSS X30Y65VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X30Y80VDD X30Y70VDD X30Y75VDD 25mOhm
L_X30Y70VDD_X30Y80VDD X30Y75VDD X30Y80VDD 2.91e-06nH
R_X30Y70VSS_X30Y80VSS X30Y70VSS X30Y75VSS 25mOhm
L_X30Y70VSS_X30Y80VSS X30Y75VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X30Y90VDD X30Y80VDD X30Y85VDD 25mOhm
L_X30Y80VDD_X30Y90VDD X30Y85VDD X30Y90VDD 2.91e-06nH
R_X30Y80VSS_X30Y90VSS X30Y80VSS X30Y85VSS 25mOhm
L_X30Y80VSS_X30Y90VSS X30Y85VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X30Y100VDD X30Y90VDD X30Y95VDD 25mOhm
L_X30Y90VDD_X30Y100VDD X30Y95VDD X30Y100VDD 2.91e-06nH
R_X30Y90VSS_X30Y100VSS X30Y90VSS X30Y95VSS 25mOhm
L_X30Y90VSS_X30Y100VSS X30Y95VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X30Y110VDD X30Y100VDD X30Y105VDD 25mOhm
L_X30Y100VDD_X30Y110VDD X30Y105VDD X30Y110VDD 2.91e-06nH
R_X30Y100VSS_X30Y110VSS X30Y100VSS X30Y105VSS 25mOhm
L_X30Y100VSS_X30Y110VSS X30Y105VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X30Y120VDD X30Y110VDD X30Y115VDD 25mOhm
L_X30Y110VDD_X30Y120VDD X30Y115VDD X30Y120VDD 2.91e-06nH
R_X30Y110VSS_X30Y120VSS X30Y110VSS X30Y115VSS 25mOhm
L_X30Y110VSS_X30Y120VSS X30Y115VSS X30Y120VSS 2.91e-06nH
R_X40Y10VDD_X40Y20VDD X40Y10VDD X40Y15VDD 25mOhm
L_X40Y10VDD_X40Y20VDD X40Y15VDD X40Y20VDD 2.91e-06nH
R_X40Y10VSS_X40Y20VSS X40Y10VSS X40Y15VSS 25mOhm
L_X40Y10VSS_X40Y20VSS X40Y15VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X40Y30VDD X40Y20VDD X40Y25VDD 25mOhm
L_X40Y20VDD_X40Y30VDD X40Y25VDD X40Y30VDD 2.91e-06nH
R_X40Y20VSS_X40Y30VSS X40Y20VSS X40Y25VSS 25mOhm
L_X40Y20VSS_X40Y30VSS X40Y25VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X40Y40VDD X40Y30VDD X40Y35VDD 25mOhm
L_X40Y30VDD_X40Y40VDD X40Y35VDD X40Y40VDD 2.91e-06nH
R_X40Y30VSS_X40Y40VSS X40Y30VSS X40Y35VSS 25mOhm
L_X40Y30VSS_X40Y40VSS X40Y35VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X40Y50VDD X40Y40VDD X40Y45VDD 25mOhm
L_X40Y40VDD_X40Y50VDD X40Y45VDD X40Y50VDD 2.91e-06nH
R_X40Y40VSS_X40Y50VSS X40Y40VSS X40Y45VSS 25mOhm
L_X40Y40VSS_X40Y50VSS X40Y45VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X40Y60VDD X40Y50VDD X40Y55VDD 25mOhm
L_X40Y50VDD_X40Y60VDD X40Y55VDD X40Y60VDD 2.91e-06nH
R_X40Y50VSS_X40Y60VSS X40Y50VSS X40Y55VSS 25mOhm
L_X40Y50VSS_X40Y60VSS X40Y55VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X40Y70VDD X40Y60VDD X40Y65VDD 25mOhm
L_X40Y60VDD_X40Y70VDD X40Y65VDD X40Y70VDD 2.91e-06nH
R_X40Y60VSS_X40Y70VSS X40Y60VSS X40Y65VSS 25mOhm
L_X40Y60VSS_X40Y70VSS X40Y65VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X40Y80VDD X40Y70VDD X40Y75VDD 25mOhm
L_X40Y70VDD_X40Y80VDD X40Y75VDD X40Y80VDD 2.91e-06nH
R_X40Y70VSS_X40Y80VSS X40Y70VSS X40Y75VSS 25mOhm
L_X40Y70VSS_X40Y80VSS X40Y75VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X40Y90VDD X40Y80VDD X40Y85VDD 25mOhm
L_X40Y80VDD_X40Y90VDD X40Y85VDD X40Y90VDD 2.91e-06nH
R_X40Y80VSS_X40Y90VSS X40Y80VSS X40Y85VSS 25mOhm
L_X40Y80VSS_X40Y90VSS X40Y85VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X40Y100VDD X40Y90VDD X40Y95VDD 25mOhm
L_X40Y90VDD_X40Y100VDD X40Y95VDD X40Y100VDD 2.91e-06nH
R_X40Y90VSS_X40Y100VSS X40Y90VSS X40Y95VSS 25mOhm
L_X40Y90VSS_X40Y100VSS X40Y95VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X40Y110VDD X40Y100VDD X40Y105VDD 25mOhm
L_X40Y100VDD_X40Y110VDD X40Y105VDD X40Y110VDD 2.91e-06nH
R_X40Y100VSS_X40Y110VSS X40Y100VSS X40Y105VSS 25mOhm
L_X40Y100VSS_X40Y110VSS X40Y105VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X40Y120VDD X40Y110VDD X40Y115VDD 25mOhm
L_X40Y110VDD_X40Y120VDD X40Y115VDD X40Y120VDD 2.91e-06nH
R_X40Y110VSS_X40Y120VSS X40Y110VSS X40Y115VSS 25mOhm
L_X40Y110VSS_X40Y120VSS X40Y115VSS X40Y120VSS 2.91e-06nH
R_X50Y10VDD_X50Y20VDD X50Y10VDD X50Y15VDD 25mOhm
L_X50Y10VDD_X50Y20VDD X50Y15VDD X50Y20VDD 2.91e-06nH
R_X50Y10VSS_X50Y20VSS X50Y10VSS X50Y15VSS 25mOhm
L_X50Y10VSS_X50Y20VSS X50Y15VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X50Y30VDD X50Y20VDD X50Y25VDD 25mOhm
L_X50Y20VDD_X50Y30VDD X50Y25VDD X50Y30VDD 2.91e-06nH
R_X50Y20VSS_X50Y30VSS X50Y20VSS X50Y25VSS 25mOhm
L_X50Y20VSS_X50Y30VSS X50Y25VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X50Y40VDD X50Y30VDD X50Y35VDD 25mOhm
L_X50Y30VDD_X50Y40VDD X50Y35VDD X50Y40VDD 2.91e-06nH
R_X50Y30VSS_X50Y40VSS X50Y30VSS X50Y35VSS 25mOhm
L_X50Y30VSS_X50Y40VSS X50Y35VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X50Y50VDD X50Y40VDD X50Y45VDD 25mOhm
L_X50Y40VDD_X50Y50VDD X50Y45VDD X50Y50VDD 2.91e-06nH
R_X50Y40VSS_X50Y50VSS X50Y40VSS X50Y45VSS 25mOhm
L_X50Y40VSS_X50Y50VSS X50Y45VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X50Y60VDD X50Y50VDD X50Y55VDD 25mOhm
L_X50Y50VDD_X50Y60VDD X50Y55VDD X50Y60VDD 2.91e-06nH
R_X50Y50VSS_X50Y60VSS X50Y50VSS X50Y55VSS 25mOhm
L_X50Y50VSS_X50Y60VSS X50Y55VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X50Y70VDD X50Y60VDD X50Y65VDD 25mOhm
L_X50Y60VDD_X50Y70VDD X50Y65VDD X50Y70VDD 2.91e-06nH
R_X50Y60VSS_X50Y70VSS X50Y60VSS X50Y65VSS 25mOhm
L_X50Y60VSS_X50Y70VSS X50Y65VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X50Y80VDD X50Y70VDD X50Y75VDD 25mOhm
L_X50Y70VDD_X50Y80VDD X50Y75VDD X50Y80VDD 2.91e-06nH
R_X50Y70VSS_X50Y80VSS X50Y70VSS X50Y75VSS 25mOhm
L_X50Y70VSS_X50Y80VSS X50Y75VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X50Y90VDD X50Y80VDD X50Y85VDD 25mOhm
L_X50Y80VDD_X50Y90VDD X50Y85VDD X50Y90VDD 2.91e-06nH
R_X50Y80VSS_X50Y90VSS X50Y80VSS X50Y85VSS 25mOhm
L_X50Y80VSS_X50Y90VSS X50Y85VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X50Y100VDD X50Y90VDD X50Y95VDD 25mOhm
L_X50Y90VDD_X50Y100VDD X50Y95VDD X50Y100VDD 2.91e-06nH
R_X50Y90VSS_X50Y100VSS X50Y90VSS X50Y95VSS 25mOhm
L_X50Y90VSS_X50Y100VSS X50Y95VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X50Y110VDD X50Y100VDD X50Y105VDD 25mOhm
L_X50Y100VDD_X50Y110VDD X50Y105VDD X50Y110VDD 2.91e-06nH
R_X50Y100VSS_X50Y110VSS X50Y100VSS X50Y105VSS 25mOhm
L_X50Y100VSS_X50Y110VSS X50Y105VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X50Y120VDD X50Y110VDD X50Y115VDD 25mOhm
L_X50Y110VDD_X50Y120VDD X50Y115VDD X50Y120VDD 2.91e-06nH
R_X50Y110VSS_X50Y120VSS X50Y110VSS X50Y115VSS 25mOhm
L_X50Y110VSS_X50Y120VSS X50Y115VSS X50Y120VSS 2.91e-06nH
R_X60Y10VDD_X60Y20VDD X60Y10VDD X60Y15VDD 25mOhm
L_X60Y10VDD_X60Y20VDD X60Y15VDD X60Y20VDD 2.91e-06nH
R_X60Y10VSS_X60Y20VSS X60Y10VSS X60Y15VSS 25mOhm
L_X60Y10VSS_X60Y20VSS X60Y15VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X60Y30VDD X60Y20VDD X60Y25VDD 25mOhm
L_X60Y20VDD_X60Y30VDD X60Y25VDD X60Y30VDD 2.91e-06nH
R_X60Y20VSS_X60Y30VSS X60Y20VSS X60Y25VSS 25mOhm
L_X60Y20VSS_X60Y30VSS X60Y25VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X60Y40VDD X60Y30VDD X60Y35VDD 25mOhm
L_X60Y30VDD_X60Y40VDD X60Y35VDD X60Y40VDD 2.91e-06nH
R_X60Y30VSS_X60Y40VSS X60Y30VSS X60Y35VSS 25mOhm
L_X60Y30VSS_X60Y40VSS X60Y35VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X60Y50VDD X60Y40VDD X60Y45VDD 25mOhm
L_X60Y40VDD_X60Y50VDD X60Y45VDD X60Y50VDD 2.91e-06nH
R_X60Y40VSS_X60Y50VSS X60Y40VSS X60Y45VSS 25mOhm
L_X60Y40VSS_X60Y50VSS X60Y45VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X60Y60VDD X60Y50VDD X60Y55VDD 25mOhm
L_X60Y50VDD_X60Y60VDD X60Y55VDD X60Y60VDD 2.91e-06nH
R_X60Y50VSS_X60Y60VSS X60Y50VSS X60Y55VSS 25mOhm
L_X60Y50VSS_X60Y60VSS X60Y55VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X60Y70VDD X60Y60VDD X60Y65VDD 25mOhm
L_X60Y60VDD_X60Y70VDD X60Y65VDD X60Y70VDD 2.91e-06nH
R_X60Y60VSS_X60Y70VSS X60Y60VSS X60Y65VSS 25mOhm
L_X60Y60VSS_X60Y70VSS X60Y65VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X60Y80VDD X60Y70VDD X60Y75VDD 25mOhm
L_X60Y70VDD_X60Y80VDD X60Y75VDD X60Y80VDD 2.91e-06nH
R_X60Y70VSS_X60Y80VSS X60Y70VSS X60Y75VSS 25mOhm
L_X60Y70VSS_X60Y80VSS X60Y75VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X60Y90VDD X60Y80VDD X60Y85VDD 25mOhm
L_X60Y80VDD_X60Y90VDD X60Y85VDD X60Y90VDD 2.91e-06nH
R_X60Y80VSS_X60Y90VSS X60Y80VSS X60Y85VSS 25mOhm
L_X60Y80VSS_X60Y90VSS X60Y85VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X60Y100VDD X60Y90VDD X60Y95VDD 25mOhm
L_X60Y90VDD_X60Y100VDD X60Y95VDD X60Y100VDD 2.91e-06nH
R_X60Y90VSS_X60Y100VSS X60Y90VSS X60Y95VSS 25mOhm
L_X60Y90VSS_X60Y100VSS X60Y95VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X60Y110VDD X60Y100VDD X60Y105VDD 25mOhm
L_X60Y100VDD_X60Y110VDD X60Y105VDD X60Y110VDD 2.91e-06nH
R_X60Y100VSS_X60Y110VSS X60Y100VSS X60Y105VSS 25mOhm
L_X60Y100VSS_X60Y110VSS X60Y105VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X60Y120VDD X60Y110VDD X60Y115VDD 25mOhm
L_X60Y110VDD_X60Y120VDD X60Y115VDD X60Y120VDD 2.91e-06nH
R_X60Y110VSS_X60Y120VSS X60Y110VSS X60Y115VSS 25mOhm
L_X60Y110VSS_X60Y120VSS X60Y115VSS X60Y120VSS 2.91e-06nH
R_X70Y10VDD_X70Y20VDD X70Y10VDD X70Y15VDD 25mOhm
L_X70Y10VDD_X70Y20VDD X70Y15VDD X70Y20VDD 2.91e-06nH
R_X70Y10VSS_X70Y20VSS X70Y10VSS X70Y15VSS 25mOhm
L_X70Y10VSS_X70Y20VSS X70Y15VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X70Y30VDD X70Y20VDD X70Y25VDD 25mOhm
L_X70Y20VDD_X70Y30VDD X70Y25VDD X70Y30VDD 2.91e-06nH
R_X70Y20VSS_X70Y30VSS X70Y20VSS X70Y25VSS 25mOhm
L_X70Y20VSS_X70Y30VSS X70Y25VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X70Y40VDD X70Y30VDD X70Y35VDD 25mOhm
L_X70Y30VDD_X70Y40VDD X70Y35VDD X70Y40VDD 2.91e-06nH
R_X70Y30VSS_X70Y40VSS X70Y30VSS X70Y35VSS 25mOhm
L_X70Y30VSS_X70Y40VSS X70Y35VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X70Y50VDD X70Y40VDD X70Y45VDD 25mOhm
L_X70Y40VDD_X70Y50VDD X70Y45VDD X70Y50VDD 2.91e-06nH
R_X70Y40VSS_X70Y50VSS X70Y40VSS X70Y45VSS 25mOhm
L_X70Y40VSS_X70Y50VSS X70Y45VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X70Y60VDD X70Y50VDD X70Y55VDD 25mOhm
L_X70Y50VDD_X70Y60VDD X70Y55VDD X70Y60VDD 2.91e-06nH
R_X70Y50VSS_X70Y60VSS X70Y50VSS X70Y55VSS 25mOhm
L_X70Y50VSS_X70Y60VSS X70Y55VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X70Y70VDD X70Y60VDD X70Y65VDD 25mOhm
L_X70Y60VDD_X70Y70VDD X70Y65VDD X70Y70VDD 2.91e-06nH
R_X70Y60VSS_X70Y70VSS X70Y60VSS X70Y65VSS 25mOhm
L_X70Y60VSS_X70Y70VSS X70Y65VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X70Y80VDD X70Y70VDD X70Y75VDD 25mOhm
L_X70Y70VDD_X70Y80VDD X70Y75VDD X70Y80VDD 2.91e-06nH
R_X70Y70VSS_X70Y80VSS X70Y70VSS X70Y75VSS 25mOhm
L_X70Y70VSS_X70Y80VSS X70Y75VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X70Y90VDD X70Y80VDD X70Y85VDD 25mOhm
L_X70Y80VDD_X70Y90VDD X70Y85VDD X70Y90VDD 2.91e-06nH
R_X70Y80VSS_X70Y90VSS X70Y80VSS X70Y85VSS 25mOhm
L_X70Y80VSS_X70Y90VSS X70Y85VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X70Y100VDD X70Y90VDD X70Y95VDD 25mOhm
L_X70Y90VDD_X70Y100VDD X70Y95VDD X70Y100VDD 2.91e-06nH
R_X70Y90VSS_X70Y100VSS X70Y90VSS X70Y95VSS 25mOhm
L_X70Y90VSS_X70Y100VSS X70Y95VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X70Y110VDD X70Y100VDD X70Y105VDD 25mOhm
L_X70Y100VDD_X70Y110VDD X70Y105VDD X70Y110VDD 2.91e-06nH
R_X70Y100VSS_X70Y110VSS X70Y100VSS X70Y105VSS 25mOhm
L_X70Y100VSS_X70Y110VSS X70Y105VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X70Y120VDD X70Y110VDD X70Y115VDD 25mOhm
L_X70Y110VDD_X70Y120VDD X70Y115VDD X70Y120VDD 2.91e-06nH
R_X70Y110VSS_X70Y120VSS X70Y110VSS X70Y115VSS 25mOhm
L_X70Y110VSS_X70Y120VSS X70Y115VSS X70Y120VSS 2.91e-06nH
R_X80Y10VDD_X80Y20VDD X80Y10VDD X80Y15VDD 25mOhm
L_X80Y10VDD_X80Y20VDD X80Y15VDD X80Y20VDD 2.91e-06nH
R_X80Y10VSS_X80Y20VSS X80Y10VSS X80Y15VSS 25mOhm
L_X80Y10VSS_X80Y20VSS X80Y15VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X80Y30VDD X80Y20VDD X80Y25VDD 25mOhm
L_X80Y20VDD_X80Y30VDD X80Y25VDD X80Y30VDD 2.91e-06nH
R_X80Y20VSS_X80Y30VSS X80Y20VSS X80Y25VSS 25mOhm
L_X80Y20VSS_X80Y30VSS X80Y25VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X80Y40VDD X80Y30VDD X80Y35VDD 25mOhm
L_X80Y30VDD_X80Y40VDD X80Y35VDD X80Y40VDD 2.91e-06nH
R_X80Y30VSS_X80Y40VSS X80Y30VSS X80Y35VSS 25mOhm
L_X80Y30VSS_X80Y40VSS X80Y35VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X80Y50VDD X80Y40VDD X80Y45VDD 25mOhm
L_X80Y40VDD_X80Y50VDD X80Y45VDD X80Y50VDD 2.91e-06nH
R_X80Y40VSS_X80Y50VSS X80Y40VSS X80Y45VSS 25mOhm
L_X80Y40VSS_X80Y50VSS X80Y45VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X80Y60VDD X80Y50VDD X80Y55VDD 25mOhm
L_X80Y50VDD_X80Y60VDD X80Y55VDD X80Y60VDD 2.91e-06nH
R_X80Y50VSS_X80Y60VSS X80Y50VSS X80Y55VSS 25mOhm
L_X80Y50VSS_X80Y60VSS X80Y55VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X80Y70VDD X80Y60VDD X80Y65VDD 25mOhm
L_X80Y60VDD_X80Y70VDD X80Y65VDD X80Y70VDD 2.91e-06nH
R_X80Y60VSS_X80Y70VSS X80Y60VSS X80Y65VSS 25mOhm
L_X80Y60VSS_X80Y70VSS X80Y65VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X80Y80VDD X80Y70VDD X80Y75VDD 25mOhm
L_X80Y70VDD_X80Y80VDD X80Y75VDD X80Y80VDD 2.91e-06nH
R_X80Y70VSS_X80Y80VSS X80Y70VSS X80Y75VSS 25mOhm
L_X80Y70VSS_X80Y80VSS X80Y75VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X80Y90VDD X80Y80VDD X80Y85VDD 25mOhm
L_X80Y80VDD_X80Y90VDD X80Y85VDD X80Y90VDD 2.91e-06nH
R_X80Y80VSS_X80Y90VSS X80Y80VSS X80Y85VSS 25mOhm
L_X80Y80VSS_X80Y90VSS X80Y85VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X80Y100VDD X80Y90VDD X80Y95VDD 25mOhm
L_X80Y90VDD_X80Y100VDD X80Y95VDD X80Y100VDD 2.91e-06nH
R_X80Y90VSS_X80Y100VSS X80Y90VSS X80Y95VSS 25mOhm
L_X80Y90VSS_X80Y100VSS X80Y95VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X80Y110VDD X80Y100VDD X80Y105VDD 25mOhm
L_X80Y100VDD_X80Y110VDD X80Y105VDD X80Y110VDD 2.91e-06nH
R_X80Y100VSS_X80Y110VSS X80Y100VSS X80Y105VSS 25mOhm
L_X80Y100VSS_X80Y110VSS X80Y105VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X80Y120VDD X80Y110VDD X80Y115VDD 25mOhm
L_X80Y110VDD_X80Y120VDD X80Y115VDD X80Y120VDD 2.91e-06nH
R_X80Y110VSS_X80Y120VSS X80Y110VSS X80Y115VSS 25mOhm
L_X80Y110VSS_X80Y120VSS X80Y115VSS X80Y120VSS 2.91e-06nH
R_X90Y10VDD_X90Y20VDD X90Y10VDD X90Y15VDD 25mOhm
L_X90Y10VDD_X90Y20VDD X90Y15VDD X90Y20VDD 2.91e-06nH
R_X90Y10VSS_X90Y20VSS X90Y10VSS X90Y15VSS 25mOhm
L_X90Y10VSS_X90Y20VSS X90Y15VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X90Y30VDD X90Y20VDD X90Y25VDD 25mOhm
L_X90Y20VDD_X90Y30VDD X90Y25VDD X90Y30VDD 2.91e-06nH
R_X90Y20VSS_X90Y30VSS X90Y20VSS X90Y25VSS 25mOhm
L_X90Y20VSS_X90Y30VSS X90Y25VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X90Y40VDD X90Y30VDD X90Y35VDD 25mOhm
L_X90Y30VDD_X90Y40VDD X90Y35VDD X90Y40VDD 2.91e-06nH
R_X90Y30VSS_X90Y40VSS X90Y30VSS X90Y35VSS 25mOhm
L_X90Y30VSS_X90Y40VSS X90Y35VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X90Y50VDD X90Y40VDD X90Y45VDD 25mOhm
L_X90Y40VDD_X90Y50VDD X90Y45VDD X90Y50VDD 2.91e-06nH
R_X90Y40VSS_X90Y50VSS X90Y40VSS X90Y45VSS 25mOhm
L_X90Y40VSS_X90Y50VSS X90Y45VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X90Y60VDD X90Y50VDD X90Y55VDD 25mOhm
L_X90Y50VDD_X90Y60VDD X90Y55VDD X90Y60VDD 2.91e-06nH
R_X90Y50VSS_X90Y60VSS X90Y50VSS X90Y55VSS 25mOhm
L_X90Y50VSS_X90Y60VSS X90Y55VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X90Y70VDD X90Y60VDD X90Y65VDD 25mOhm
L_X90Y60VDD_X90Y70VDD X90Y65VDD X90Y70VDD 2.91e-06nH
R_X90Y60VSS_X90Y70VSS X90Y60VSS X90Y65VSS 25mOhm
L_X90Y60VSS_X90Y70VSS X90Y65VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X90Y80VDD X90Y70VDD X90Y75VDD 25mOhm
L_X90Y70VDD_X90Y80VDD X90Y75VDD X90Y80VDD 2.91e-06nH
R_X90Y70VSS_X90Y80VSS X90Y70VSS X90Y75VSS 25mOhm
L_X90Y70VSS_X90Y80VSS X90Y75VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X90Y90VDD X90Y80VDD X90Y85VDD 25mOhm
L_X90Y80VDD_X90Y90VDD X90Y85VDD X90Y90VDD 2.91e-06nH
R_X90Y80VSS_X90Y90VSS X90Y80VSS X90Y85VSS 25mOhm
L_X90Y80VSS_X90Y90VSS X90Y85VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X90Y100VDD X90Y90VDD X90Y95VDD 25mOhm
L_X90Y90VDD_X90Y100VDD X90Y95VDD X90Y100VDD 2.91e-06nH
R_X90Y90VSS_X90Y100VSS X90Y90VSS X90Y95VSS 25mOhm
L_X90Y90VSS_X90Y100VSS X90Y95VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X90Y110VDD X90Y100VDD X90Y105VDD 25mOhm
L_X90Y100VDD_X90Y110VDD X90Y105VDD X90Y110VDD 2.91e-06nH
R_X90Y100VSS_X90Y110VSS X90Y100VSS X90Y105VSS 25mOhm
L_X90Y100VSS_X90Y110VSS X90Y105VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X90Y120VDD X90Y110VDD X90Y115VDD 25mOhm
L_X90Y110VDD_X90Y120VDD X90Y115VDD X90Y120VDD 2.91e-06nH
R_X90Y110VSS_X90Y120VSS X90Y110VSS X90Y115VSS 25mOhm
L_X90Y110VSS_X90Y120VSS X90Y115VSS X90Y120VSS 2.91e-06nH
R_X100Y10VDD_X100Y20VDD X100Y10VDD X100Y15VDD 25mOhm
L_X100Y10VDD_X100Y20VDD X100Y15VDD X100Y20VDD 2.91e-06nH
R_X100Y10VSS_X100Y20VSS X100Y10VSS X100Y15VSS 25mOhm
L_X100Y10VSS_X100Y20VSS X100Y15VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X100Y30VDD X100Y20VDD X100Y25VDD 25mOhm
L_X100Y20VDD_X100Y30VDD X100Y25VDD X100Y30VDD 2.91e-06nH
R_X100Y20VSS_X100Y30VSS X100Y20VSS X100Y25VSS 25mOhm
L_X100Y20VSS_X100Y30VSS X100Y25VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X100Y40VDD X100Y30VDD X100Y35VDD 25mOhm
L_X100Y30VDD_X100Y40VDD X100Y35VDD X100Y40VDD 2.91e-06nH
R_X100Y30VSS_X100Y40VSS X100Y30VSS X100Y35VSS 25mOhm
L_X100Y30VSS_X100Y40VSS X100Y35VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X100Y50VDD X100Y40VDD X100Y45VDD 25mOhm
L_X100Y40VDD_X100Y50VDD X100Y45VDD X100Y50VDD 2.91e-06nH
R_X100Y40VSS_X100Y50VSS X100Y40VSS X100Y45VSS 25mOhm
L_X100Y40VSS_X100Y50VSS X100Y45VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X100Y60VDD X100Y50VDD X100Y55VDD 25mOhm
L_X100Y50VDD_X100Y60VDD X100Y55VDD X100Y60VDD 2.91e-06nH
R_X100Y50VSS_X100Y60VSS X100Y50VSS X100Y55VSS 25mOhm
L_X100Y50VSS_X100Y60VSS X100Y55VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X100Y70VDD X100Y60VDD X100Y65VDD 25mOhm
L_X100Y60VDD_X100Y70VDD X100Y65VDD X100Y70VDD 2.91e-06nH
R_X100Y60VSS_X100Y70VSS X100Y60VSS X100Y65VSS 25mOhm
L_X100Y60VSS_X100Y70VSS X100Y65VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X100Y80VDD X100Y70VDD X100Y75VDD 25mOhm
L_X100Y70VDD_X100Y80VDD X100Y75VDD X100Y80VDD 2.91e-06nH
R_X100Y70VSS_X100Y80VSS X100Y70VSS X100Y75VSS 25mOhm
L_X100Y70VSS_X100Y80VSS X100Y75VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X100Y90VDD X100Y80VDD X100Y85VDD 25mOhm
L_X100Y80VDD_X100Y90VDD X100Y85VDD X100Y90VDD 2.91e-06nH
R_X100Y80VSS_X100Y90VSS X100Y80VSS X100Y85VSS 25mOhm
L_X100Y80VSS_X100Y90VSS X100Y85VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X100Y100VDD X100Y90VDD X100Y95VDD 25mOhm
L_X100Y90VDD_X100Y100VDD X100Y95VDD X100Y100VDD 2.91e-06nH
R_X100Y90VSS_X100Y100VSS X100Y90VSS X100Y95VSS 25mOhm
L_X100Y90VSS_X100Y100VSS X100Y95VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X100Y110VDD X100Y100VDD X100Y105VDD 25mOhm
L_X100Y100VDD_X100Y110VDD X100Y105VDD X100Y110VDD 2.91e-06nH
R_X100Y100VSS_X100Y110VSS X100Y100VSS X100Y105VSS 25mOhm
L_X100Y100VSS_X100Y110VSS X100Y105VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X100Y120VDD X100Y110VDD X100Y115VDD 25mOhm
L_X100Y110VDD_X100Y120VDD X100Y115VDD X100Y120VDD 2.91e-06nH
R_X100Y110VSS_X100Y120VSS X100Y110VSS X100Y115VSS 25mOhm
L_X100Y110VSS_X100Y120VSS X100Y115VSS X100Y120VSS 2.91e-06nH
R_X110Y10VDD_X110Y20VDD X110Y10VDD X110Y15VDD 25mOhm
L_X110Y10VDD_X110Y20VDD X110Y15VDD X110Y20VDD 2.91e-06nH
R_X110Y10VSS_X110Y20VSS X110Y10VSS X110Y15VSS 25mOhm
L_X110Y10VSS_X110Y20VSS X110Y15VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X110Y30VDD X110Y20VDD X110Y25VDD 25mOhm
L_X110Y20VDD_X110Y30VDD X110Y25VDD X110Y30VDD 2.91e-06nH
R_X110Y20VSS_X110Y30VSS X110Y20VSS X110Y25VSS 25mOhm
L_X110Y20VSS_X110Y30VSS X110Y25VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X110Y40VDD X110Y30VDD X110Y35VDD 25mOhm
L_X110Y30VDD_X110Y40VDD X110Y35VDD X110Y40VDD 2.91e-06nH
R_X110Y30VSS_X110Y40VSS X110Y30VSS X110Y35VSS 25mOhm
L_X110Y30VSS_X110Y40VSS X110Y35VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X110Y50VDD X110Y40VDD X110Y45VDD 25mOhm
L_X110Y40VDD_X110Y50VDD X110Y45VDD X110Y50VDD 2.91e-06nH
R_X110Y40VSS_X110Y50VSS X110Y40VSS X110Y45VSS 25mOhm
L_X110Y40VSS_X110Y50VSS X110Y45VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X110Y60VDD X110Y50VDD X110Y55VDD 25mOhm
L_X110Y50VDD_X110Y60VDD X110Y55VDD X110Y60VDD 2.91e-06nH
R_X110Y50VSS_X110Y60VSS X110Y50VSS X110Y55VSS 25mOhm
L_X110Y50VSS_X110Y60VSS X110Y55VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X110Y70VDD X110Y60VDD X110Y65VDD 25mOhm
L_X110Y60VDD_X110Y70VDD X110Y65VDD X110Y70VDD 2.91e-06nH
R_X110Y60VSS_X110Y70VSS X110Y60VSS X110Y65VSS 25mOhm
L_X110Y60VSS_X110Y70VSS X110Y65VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X110Y80VDD X110Y70VDD X110Y75VDD 25mOhm
L_X110Y70VDD_X110Y80VDD X110Y75VDD X110Y80VDD 2.91e-06nH
R_X110Y70VSS_X110Y80VSS X110Y70VSS X110Y75VSS 25mOhm
L_X110Y70VSS_X110Y80VSS X110Y75VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X110Y90VDD X110Y80VDD X110Y85VDD 25mOhm
L_X110Y80VDD_X110Y90VDD X110Y85VDD X110Y90VDD 2.91e-06nH
R_X110Y80VSS_X110Y90VSS X110Y80VSS X110Y85VSS 25mOhm
L_X110Y80VSS_X110Y90VSS X110Y85VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X110Y100VDD X110Y90VDD X110Y95VDD 25mOhm
L_X110Y90VDD_X110Y100VDD X110Y95VDD X110Y100VDD 2.91e-06nH
R_X110Y90VSS_X110Y100VSS X110Y90VSS X110Y95VSS 25mOhm
L_X110Y90VSS_X110Y100VSS X110Y95VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X110Y110VDD X110Y100VDD X110Y105VDD 25mOhm
L_X110Y100VDD_X110Y110VDD X110Y105VDD X110Y110VDD 2.91e-06nH
R_X110Y100VSS_X110Y110VSS X110Y100VSS X110Y105VSS 25mOhm
L_X110Y100VSS_X110Y110VSS X110Y105VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X110Y120VDD X110Y110VDD X110Y115VDD 25mOhm
L_X110Y110VDD_X110Y120VDD X110Y115VDD X110Y120VDD 2.91e-06nH
R_X110Y110VSS_X110Y120VSS X110Y110VSS X110Y115VSS 25mOhm
L_X110Y110VSS_X110Y120VSS X110Y115VSS X110Y120VSS 2.91e-06nH
R_X120Y10VDD_X120Y20VDD X120Y10VDD X120Y15VDD 25mOhm
L_X120Y10VDD_X120Y20VDD X120Y15VDD X120Y20VDD 2.91e-06nH
R_X120Y10VSS_X120Y20VSS X120Y10VSS X120Y15VSS 25mOhm
L_X120Y10VSS_X120Y20VSS X120Y15VSS X120Y20VSS 2.91e-06nH
R_X120Y20VDD_X120Y30VDD X120Y20VDD X120Y25VDD 25mOhm
L_X120Y20VDD_X120Y30VDD X120Y25VDD X120Y30VDD 2.91e-06nH
R_X120Y20VSS_X120Y30VSS X120Y20VSS X120Y25VSS 25mOhm
L_X120Y20VSS_X120Y30VSS X120Y25VSS X120Y30VSS 2.91e-06nH
R_X120Y30VDD_X120Y40VDD X120Y30VDD X120Y35VDD 25mOhm
L_X120Y30VDD_X120Y40VDD X120Y35VDD X120Y40VDD 2.91e-06nH
R_X120Y30VSS_X120Y40VSS X120Y30VSS X120Y35VSS 25mOhm
L_X120Y30VSS_X120Y40VSS X120Y35VSS X120Y40VSS 2.91e-06nH
R_X120Y40VDD_X120Y50VDD X120Y40VDD X120Y45VDD 25mOhm
L_X120Y40VDD_X120Y50VDD X120Y45VDD X120Y50VDD 2.91e-06nH
R_X120Y40VSS_X120Y50VSS X120Y40VSS X120Y45VSS 25mOhm
L_X120Y40VSS_X120Y50VSS X120Y45VSS X120Y50VSS 2.91e-06nH
R_X120Y50VDD_X120Y60VDD X120Y50VDD X120Y55VDD 25mOhm
L_X120Y50VDD_X120Y60VDD X120Y55VDD X120Y60VDD 2.91e-06nH
R_X120Y50VSS_X120Y60VSS X120Y50VSS X120Y55VSS 25mOhm
L_X120Y50VSS_X120Y60VSS X120Y55VSS X120Y60VSS 2.91e-06nH
R_X120Y60VDD_X120Y70VDD X120Y60VDD X120Y65VDD 25mOhm
L_X120Y60VDD_X120Y70VDD X120Y65VDD X120Y70VDD 2.91e-06nH
R_X120Y60VSS_X120Y70VSS X120Y60VSS X120Y65VSS 25mOhm
L_X120Y60VSS_X120Y70VSS X120Y65VSS X120Y70VSS 2.91e-06nH
R_X120Y70VDD_X120Y80VDD X120Y70VDD X120Y75VDD 25mOhm
L_X120Y70VDD_X120Y80VDD X120Y75VDD X120Y80VDD 2.91e-06nH
R_X120Y70VSS_X120Y80VSS X120Y70VSS X120Y75VSS 25mOhm
L_X120Y70VSS_X120Y80VSS X120Y75VSS X120Y80VSS 2.91e-06nH
R_X120Y80VDD_X120Y90VDD X120Y80VDD X120Y85VDD 25mOhm
L_X120Y80VDD_X120Y90VDD X120Y85VDD X120Y90VDD 2.91e-06nH
R_X120Y80VSS_X120Y90VSS X120Y80VSS X120Y85VSS 25mOhm
L_X120Y80VSS_X120Y90VSS X120Y85VSS X120Y90VSS 2.91e-06nH
R_X120Y90VDD_X120Y100VDD X120Y90VDD X120Y95VDD 25mOhm
L_X120Y90VDD_X120Y100VDD X120Y95VDD X120Y100VDD 2.91e-06nH
R_X120Y90VSS_X120Y100VSS X120Y90VSS X120Y95VSS 25mOhm
L_X120Y90VSS_X120Y100VSS X120Y95VSS X120Y100VSS 2.91e-06nH
R_X120Y100VDD_X120Y110VDD X120Y100VDD X120Y105VDD 25mOhm
L_X120Y100VDD_X120Y110VDD X120Y105VDD X120Y110VDD 2.91e-06nH
R_X120Y100VSS_X120Y110VSS X120Y100VSS X120Y105VSS 25mOhm
L_X120Y100VSS_X120Y110VSS X120Y105VSS X120Y110VSS 2.91e-06nH
R_X120Y110VDD_X120Y120VDD X120Y110VDD X120Y115VDD 25mOhm
L_X120Y110VDD_X120Y120VDD X120Y115VDD X120Y120VDD 2.91e-06nH
R_X120Y110VSS_X120Y120VSS X120Y110VSS X120Y115VSS 25mOhm
L_X120Y110VSS_X120Y120VSS X120Y115VSS X120Y120VSS 2.91e-06nH
C_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VSS 10nF
C_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VSS 10nF
C_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VSS 10nF
C_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VSS 10nF
C_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VSS 10nF
C_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VSS 10nF
C_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VSS 10nF
C_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VSS 10nF
C_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VSS 10nF
C_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VSS 10nF
C_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VSS 10nF
C_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VSS 10nF
C_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VSS 10nF
C_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VSS 10nF
C_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VSS 10nF
C_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VSS 10nF
C_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VSS 10nF
C_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VSS 10nF
C_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VSS 10nF
C_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VSS 10nF
C_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VSS 10nF
C_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VSS 10nF
C_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VSS 10nF
C_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VSS 10nF
C_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VSS 10nF
C_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VSS 10nF
C_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VSS 10nF
C_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VSS 10nF
C_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VSS 10nF
C_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VSS 10nF
C_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VSS 10nF
C_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VSS 10nF
C_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VSS 10nF
C_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VSS 10nF
C_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VSS 10nF
C_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VSS 10nF
C_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VSS 10nF
C_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VSS 10nF
C_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VSS 10nF
C_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VSS 10nF
C_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VSS 10nF
C_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VSS 10nF
C_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VSS 10nF
C_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VSS 10nF
C_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VSS 10nF
C_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VSS 10nF
C_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VSS 10nF
C_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VSS 10nF
C_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VSS 10nF
C_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VSS 10nF
C_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VSS 10nF
C_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VSS 10nF
C_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VSS 10nF
C_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VSS 10nF
C_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VSS 10nF
C_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VSS 10nF
C_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VSS 10nF
C_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VSS 10nF
C_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VSS 10nF
C_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VSS 10nF
C_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VSS 10nF
C_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VSS 10nF
C_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VSS 10nF
C_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VSS 10nF
C_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VSS 10nF
C_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VSS 10nF
C_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VSS 10nF
C_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VSS 10nF
C_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VSS 10nF
C_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VSS 10nF
C_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VSS 10nF
C_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VSS 10nF
C_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VSS 10nF
C_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VSS 10nF
C_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VSS 10nF
C_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VSS 10nF
C_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VSS 10nF
C_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VSS 10nF
C_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VSS 10nF
C_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VSS 10nF
C_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VSS 10nF
C_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VSS 10nF
C_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VSS 10nF
C_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VSS 10nF
C_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VSS 10nF
C_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VSS 10nF
C_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VSS 10nF
C_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VSS 10nF
C_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VSS 10nF
C_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VSS 10nF
C_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VSS 10nF
C_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VSS 10nF
C_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VSS 10nF
C_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VSS 10nF
C_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VSS 10nF
C_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VSS 10nF
C_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VSS 10nF
C_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VSS 10nF
C_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VSS 10nF
C_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VSS 10nF
C_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VSS 10nF
C_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VSS 10nF
C_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VSS 10nF
C_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VSS 10nF
C_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VSS 10nF
C_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VSS 10nF
C_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VSS 10nF
C_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VSS 10nF
C_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VSS 10nF
C_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VSS 10nF
C_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VSS 10nF
C_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VSS 10nF
C_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VSS 10nF
C_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VSS 10nF
C_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VSS 10nF
C_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VSS 10nF
C_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VSS 10nF
C_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VSS 10nF
C_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VSS 10nF
C_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VSS 10nF
C_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VSS 10nF
C_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VSS 10nF
C_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VSS 10nF
C_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VSS 10nF
C_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VSS 10nF
C_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VSS 10nF
C_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VSS 10nF
C_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VSS 10nF
C_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VSS 10nF
C_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VSS 10nF
C_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VSS 10nF
C_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VSS 10nF
C_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VSS 10nF
C_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VSS 10nF
C_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VSS 10nF
C_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VSS 10nF
C_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VSS 10nF
C_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VSS 10nF
C_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VSS 10nF
C_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VSS 10nF
C_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VSS 10nF
C_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VSS 10nF
C_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VSS 10nF
C_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VSS 10nF
I_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VDDDM 0.8 AC=1
V_X120Y120VDD_X120Y120VSS X120Y120VDDDM X120Y120VSS 0
I_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VDDDM 0.8 AC=1
V_X120Y10VDD_X120Y10VSS X120Y10VDDDM X120Y10VSS 0
I_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VDDDM 0.8 AC=1
V_X120Y20VDD_X120Y20VSS X120Y20VDDDM X120Y20VSS 0
I_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VDDDM 0.8 AC=1
V_X120Y30VDD_X120Y30VSS X120Y30VDDDM X120Y30VSS 0
I_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VDDDM 0.8 AC=1
V_X120Y40VDD_X120Y40VSS X120Y40VDDDM X120Y40VSS 0
I_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VDDDM 0.8 AC=1
V_X120Y50VDD_X120Y50VSS X120Y50VDDDM X120Y50VSS 0
I_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VDDDM 0.8 AC=1
V_X120Y60VDD_X120Y60VSS X120Y60VDDDM X120Y60VSS 0
I_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VDDDM 0.8 AC=1
V_X120Y70VDD_X120Y70VSS X120Y70VDDDM X120Y70VSS 0
I_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VDDDM 0.8 AC=1
V_X120Y80VDD_X120Y80VSS X120Y80VDDDM X120Y80VSS 0
I_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VDDDM 0.8 AC=1
V_X120Y90VDD_X120Y90VSS X120Y90VDDDM X120Y90VSS 0
I_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VDDDM 0.8 AC=1
V_X120Y100VDD_X120Y100VSS X120Y100VDDDM X120Y100VSS 0
I_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VDDDM 0.8 AC=1
V_X120Y110VDD_X120Y110VSS X120Y110VDDDM X120Y110VSS 0
I_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VDDDM 0.8 AC=1
V_X10Y120VDD_X10Y120VSS X10Y120VDDDM X10Y120VSS 0
I_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VDDDM 0.8 AC=1
V_X10Y10VDD_X10Y10VSS X10Y10VDDDM X10Y10VSS 0
I_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VDDDM 0.8 AC=1
V_X10Y20VDD_X10Y20VSS X10Y20VDDDM X10Y20VSS 0
I_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VDDDM 0.8 AC=1
V_X10Y30VDD_X10Y30VSS X10Y30VDDDM X10Y30VSS 0
I_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VDDDM 0.8 AC=1
V_X10Y40VDD_X10Y40VSS X10Y40VDDDM X10Y40VSS 0
I_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VDDDM 0.8 AC=1
V_X10Y50VDD_X10Y50VSS X10Y50VDDDM X10Y50VSS 0
I_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VDDDM 0.8 AC=1
V_X10Y60VDD_X10Y60VSS X10Y60VDDDM X10Y60VSS 0
I_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VDDDM 0.8 AC=1
V_X10Y70VDD_X10Y70VSS X10Y70VDDDM X10Y70VSS 0
I_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VDDDM 0.8 AC=1
V_X10Y80VDD_X10Y80VSS X10Y80VDDDM X10Y80VSS 0
I_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VDDDM 0.8 AC=1
V_X10Y90VDD_X10Y90VSS X10Y90VDDDM X10Y90VSS 0
I_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VDDDM 0.8 AC=1
V_X10Y100VDD_X10Y100VSS X10Y100VDDDM X10Y100VSS 0
I_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VDDDM 0.8 AC=1
V_X10Y110VDD_X10Y110VSS X10Y110VDDDM X10Y110VSS 0
I_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VDDDM 0.8 AC=1
V_X20Y120VDD_X20Y120VSS X20Y120VDDDM X20Y120VSS 0
I_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VDDDM 0.8 AC=1
V_X20Y10VDD_X20Y10VSS X20Y10VDDDM X20Y10VSS 0
I_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VDDDM 0.8 AC=1
V_X20Y20VDD_X20Y20VSS X20Y20VDDDM X20Y20VSS 0
I_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VDDDM 0.8 AC=1
V_X20Y30VDD_X20Y30VSS X20Y30VDDDM X20Y30VSS 0
I_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VDDDM 0.8 AC=1
V_X20Y40VDD_X20Y40VSS X20Y40VDDDM X20Y40VSS 0
I_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VDDDM 0.8 AC=1
V_X20Y50VDD_X20Y50VSS X20Y50VDDDM X20Y50VSS 0
I_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VDDDM 0.8 AC=1
V_X20Y60VDD_X20Y60VSS X20Y60VDDDM X20Y60VSS 0
I_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VDDDM 0.8 AC=1
V_X20Y70VDD_X20Y70VSS X20Y70VDDDM X20Y70VSS 0
I_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VDDDM 0.8 AC=1
V_X20Y80VDD_X20Y80VSS X20Y80VDDDM X20Y80VSS 0
I_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VDDDM 0.8 AC=1
V_X20Y90VDD_X20Y90VSS X20Y90VDDDM X20Y90VSS 0
I_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VDDDM 0.8 AC=1
V_X20Y100VDD_X20Y100VSS X20Y100VDDDM X20Y100VSS 0
I_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VDDDM 0.8 AC=1
V_X20Y110VDD_X20Y110VSS X20Y110VDDDM X20Y110VSS 0
I_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VDDDM 0.8 AC=1
V_X30Y120VDD_X30Y120VSS X30Y120VDDDM X30Y120VSS 0
I_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VDDDM 0.8 AC=1
V_X30Y10VDD_X30Y10VSS X30Y10VDDDM X30Y10VSS 0
I_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VDDDM 0.8 AC=1
V_X30Y20VDD_X30Y20VSS X30Y20VDDDM X30Y20VSS 0
I_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VDDDM 0.8 AC=1
V_X30Y30VDD_X30Y30VSS X30Y30VDDDM X30Y30VSS 0
I_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VDDDM 0.8 AC=1
V_X30Y40VDD_X30Y40VSS X30Y40VDDDM X30Y40VSS 0
I_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VDDDM 0.8 AC=1
V_X30Y50VDD_X30Y50VSS X30Y50VDDDM X30Y50VSS 0
I_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VDDDM 0.8 AC=1
V_X30Y60VDD_X30Y60VSS X30Y60VDDDM X30Y60VSS 0
I_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VDDDM 0.8 AC=1
V_X30Y70VDD_X30Y70VSS X30Y70VDDDM X30Y70VSS 0
I_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VDDDM 0.8 AC=1
V_X30Y80VDD_X30Y80VSS X30Y80VDDDM X30Y80VSS 0
I_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VDDDM 0.8 AC=1
V_X30Y90VDD_X30Y90VSS X30Y90VDDDM X30Y90VSS 0
I_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VDDDM 0.8 AC=1
V_X30Y100VDD_X30Y100VSS X30Y100VDDDM X30Y100VSS 0
I_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VDDDM 0.8 AC=1
V_X30Y110VDD_X30Y110VSS X30Y110VDDDM X30Y110VSS 0
I_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VDDDM 0.8 AC=1
V_X40Y120VDD_X40Y120VSS X40Y120VDDDM X40Y120VSS 0
I_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VDDDM 0.8 AC=1
V_X40Y10VDD_X40Y10VSS X40Y10VDDDM X40Y10VSS 0
I_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VDDDM 0.8 AC=1
V_X40Y20VDD_X40Y20VSS X40Y20VDDDM X40Y20VSS 0
I_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VDDDM 0.8 AC=1
V_X40Y30VDD_X40Y30VSS X40Y30VDDDM X40Y30VSS 0
I_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VDDDM 0.8 AC=1
V_X40Y40VDD_X40Y40VSS X40Y40VDDDM X40Y40VSS 0
I_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VDDDM 0.8 AC=1
V_X40Y50VDD_X40Y50VSS X40Y50VDDDM X40Y50VSS 0
I_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VDDDM 0.8 AC=1
V_X40Y60VDD_X40Y60VSS X40Y60VDDDM X40Y60VSS 0
I_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VDDDM 0.8 AC=1
V_X40Y70VDD_X40Y70VSS X40Y70VDDDM X40Y70VSS 0
I_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VDDDM 0.8 AC=1
V_X40Y80VDD_X40Y80VSS X40Y80VDDDM X40Y80VSS 0
I_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VDDDM 0.8 AC=1
V_X40Y90VDD_X40Y90VSS X40Y90VDDDM X40Y90VSS 0
I_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VDDDM 0.8 AC=1
V_X40Y100VDD_X40Y100VSS X40Y100VDDDM X40Y100VSS 0
I_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VDDDM 0.8 AC=1
V_X40Y110VDD_X40Y110VSS X40Y110VDDDM X40Y110VSS 0
I_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VDDDM 0.8 AC=1
V_X50Y120VDD_X50Y120VSS X50Y120VDDDM X50Y120VSS 0
I_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VDDDM 0.8 AC=1
V_X50Y10VDD_X50Y10VSS X50Y10VDDDM X50Y10VSS 0
I_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VDDDM 0.8 AC=1
V_X50Y20VDD_X50Y20VSS X50Y20VDDDM X50Y20VSS 0
I_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VDDDM 0.8 AC=1
V_X50Y30VDD_X50Y30VSS X50Y30VDDDM X50Y30VSS 0
I_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VDDDM 0.8 AC=1
V_X50Y40VDD_X50Y40VSS X50Y40VDDDM X50Y40VSS 0
I_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VDDDM 0.8 AC=1
V_X50Y50VDD_X50Y50VSS X50Y50VDDDM X50Y50VSS 0
I_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VDDDM 0.8 AC=1
V_X50Y60VDD_X50Y60VSS X50Y60VDDDM X50Y60VSS 0
I_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VDDDM 0.8 AC=1
V_X50Y70VDD_X50Y70VSS X50Y70VDDDM X50Y70VSS 0
I_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VDDDM 0.8 AC=1
V_X50Y80VDD_X50Y80VSS X50Y80VDDDM X50Y80VSS 0
I_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VDDDM 0.8 AC=1
V_X50Y90VDD_X50Y90VSS X50Y90VDDDM X50Y90VSS 0
I_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VDDDM 0.8 AC=1
V_X50Y100VDD_X50Y100VSS X50Y100VDDDM X50Y100VSS 0
I_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VDDDM 0.8 AC=1
V_X50Y110VDD_X50Y110VSS X50Y110VDDDM X50Y110VSS 0
I_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VDDDM 0.8 AC=1
V_X60Y120VDD_X60Y120VSS X60Y120VDDDM X60Y120VSS 0
I_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VDDDM 0.8 AC=1
V_X60Y10VDD_X60Y10VSS X60Y10VDDDM X60Y10VSS 0
I_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VDDDM 0.8 AC=1
V_X60Y20VDD_X60Y20VSS X60Y20VDDDM X60Y20VSS 0
I_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VDDDM 0.8 AC=1
V_X60Y30VDD_X60Y30VSS X60Y30VDDDM X60Y30VSS 0
I_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VDDDM 0.8 AC=1
V_X60Y40VDD_X60Y40VSS X60Y40VDDDM X60Y40VSS 0
I_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VDDDM 0.8 AC=1
V_X60Y50VDD_X60Y50VSS X60Y50VDDDM X60Y50VSS 0
I_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VDDDM 0.8 AC=1
V_X60Y60VDD_X60Y60VSS X60Y60VDDDM X60Y60VSS 0
I_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VDDDM 0.8 AC=1
V_X60Y70VDD_X60Y70VSS X60Y70VDDDM X60Y70VSS 0
I_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VDDDM 0.8 AC=1
V_X60Y80VDD_X60Y80VSS X60Y80VDDDM X60Y80VSS 0
I_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VDDDM 0.8 AC=1
V_X60Y90VDD_X60Y90VSS X60Y90VDDDM X60Y90VSS 0
I_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VDDDM 0.8 AC=1
V_X60Y100VDD_X60Y100VSS X60Y100VDDDM X60Y100VSS 0
I_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VDDDM 0.8 AC=1
V_X60Y110VDD_X60Y110VSS X60Y110VDDDM X60Y110VSS 0
I_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VDDDM 0.8 AC=1
V_X70Y120VDD_X70Y120VSS X70Y120VDDDM X70Y120VSS 0
I_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VDDDM 0.8 AC=1
V_X70Y10VDD_X70Y10VSS X70Y10VDDDM X70Y10VSS 0
I_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VDDDM 0.8 AC=1
V_X70Y20VDD_X70Y20VSS X70Y20VDDDM X70Y20VSS 0
I_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VDDDM 0.8 AC=1
V_X70Y30VDD_X70Y30VSS X70Y30VDDDM X70Y30VSS 0
I_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VDDDM 0.8 AC=1
V_X70Y40VDD_X70Y40VSS X70Y40VDDDM X70Y40VSS 0
I_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VDDDM 0.8 AC=1
V_X70Y50VDD_X70Y50VSS X70Y50VDDDM X70Y50VSS 0
I_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VDDDM 0.8 AC=1
V_X70Y60VDD_X70Y60VSS X70Y60VDDDM X70Y60VSS 0
I_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VDDDM 0.8 AC=1
V_X70Y70VDD_X70Y70VSS X70Y70VDDDM X70Y70VSS 0
I_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VDDDM 0.8 AC=1
V_X70Y80VDD_X70Y80VSS X70Y80VDDDM X70Y80VSS 0
I_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VDDDM 0.8 AC=1
V_X70Y90VDD_X70Y90VSS X70Y90VDDDM X70Y90VSS 0
I_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VDDDM 0.8 AC=1
V_X70Y100VDD_X70Y100VSS X70Y100VDDDM X70Y100VSS 0
I_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VDDDM 0.8 AC=1
V_X70Y110VDD_X70Y110VSS X70Y110VDDDM X70Y110VSS 0
I_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VDDDM 0.8 AC=1
V_X80Y120VDD_X80Y120VSS X80Y120VDDDM X80Y120VSS 0
I_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VDDDM 0.8 AC=1
V_X80Y10VDD_X80Y10VSS X80Y10VDDDM X80Y10VSS 0
I_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VDDDM 0.8 AC=1
V_X80Y20VDD_X80Y20VSS X80Y20VDDDM X80Y20VSS 0
I_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VDDDM 0.8 AC=1
V_X80Y30VDD_X80Y30VSS X80Y30VDDDM X80Y30VSS 0
I_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VDDDM 0.8 AC=1
V_X80Y40VDD_X80Y40VSS X80Y40VDDDM X80Y40VSS 0
I_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VDDDM 0.8 AC=1
V_X80Y50VDD_X80Y50VSS X80Y50VDDDM X80Y50VSS 0
I_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VDDDM 0.8 AC=1
V_X80Y60VDD_X80Y60VSS X80Y60VDDDM X80Y60VSS 0
I_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VDDDM 0.8 AC=1
V_X80Y70VDD_X80Y70VSS X80Y70VDDDM X80Y70VSS 0
I_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VDDDM 0.8 AC=1
V_X80Y80VDD_X80Y80VSS X80Y80VDDDM X80Y80VSS 0
I_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VDDDM 0.8 AC=1
V_X80Y90VDD_X80Y90VSS X80Y90VDDDM X80Y90VSS 0
I_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VDDDM 0.8 AC=1
V_X80Y100VDD_X80Y100VSS X80Y100VDDDM X80Y100VSS 0
I_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VDDDM 0.8 AC=1
V_X80Y110VDD_X80Y110VSS X80Y110VDDDM X80Y110VSS 0
I_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VDDDM 0.8 AC=1
V_X90Y120VDD_X90Y120VSS X90Y120VDDDM X90Y120VSS 0
I_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VDDDM 0.8 AC=1
V_X90Y10VDD_X90Y10VSS X90Y10VDDDM X90Y10VSS 0
I_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VDDDM 0.8 AC=1
V_X90Y20VDD_X90Y20VSS X90Y20VDDDM X90Y20VSS 0
I_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VDDDM 0.8 AC=1
V_X90Y30VDD_X90Y30VSS X90Y30VDDDM X90Y30VSS 0
I_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VDDDM 0.8 AC=1
V_X90Y40VDD_X90Y40VSS X90Y40VDDDM X90Y40VSS 0
I_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VDDDM 0.8 AC=1
V_X90Y50VDD_X90Y50VSS X90Y50VDDDM X90Y50VSS 0
I_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VDDDM 0.8 AC=1
V_X90Y60VDD_X90Y60VSS X90Y60VDDDM X90Y60VSS 0
I_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VDDDM 0.8 AC=1
V_X90Y70VDD_X90Y70VSS X90Y70VDDDM X90Y70VSS 0
I_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VDDDM 0.8 AC=1
V_X90Y80VDD_X90Y80VSS X90Y80VDDDM X90Y80VSS 0
I_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VDDDM 0.8 AC=1
V_X90Y90VDD_X90Y90VSS X90Y90VDDDM X90Y90VSS 0
I_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VDDDM 0.8 AC=1
V_X90Y100VDD_X90Y100VSS X90Y100VDDDM X90Y100VSS 0
I_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VDDDM 0.8 AC=1
V_X90Y110VDD_X90Y110VSS X90Y110VDDDM X90Y110VSS 0
I_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VDDDM 0.8 AC=1
V_X100Y120VDD_X100Y120VSS X100Y120VDDDM X100Y120VSS 0
I_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VDDDM 0.8 AC=1
V_X100Y10VDD_X100Y10VSS X100Y10VDDDM X100Y10VSS 0
I_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VDDDM 0.8 AC=1
V_X100Y20VDD_X100Y20VSS X100Y20VDDDM X100Y20VSS 0
I_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VDDDM 0.8 AC=1
V_X100Y30VDD_X100Y30VSS X100Y30VDDDM X100Y30VSS 0
I_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VDDDM 0.8 AC=1
V_X100Y40VDD_X100Y40VSS X100Y40VDDDM X100Y40VSS 0
I_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VDDDM 0.8 AC=1
V_X100Y50VDD_X100Y50VSS X100Y50VDDDM X100Y50VSS 0
I_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VDDDM 0.8 AC=1
V_X100Y60VDD_X100Y60VSS X100Y60VDDDM X100Y60VSS 0
I_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VDDDM 0.8 AC=1
V_X100Y70VDD_X100Y70VSS X100Y70VDDDM X100Y70VSS 0
I_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VDDDM 0.8 AC=1
V_X100Y80VDD_X100Y80VSS X100Y80VDDDM X100Y80VSS 0
I_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VDDDM 0.8 AC=1
V_X100Y90VDD_X100Y90VSS X100Y90VDDDM X100Y90VSS 0
I_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VDDDM 0.8 AC=1
V_X100Y100VDD_X100Y100VSS X100Y100VDDDM X100Y100VSS 0
I_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VDDDM 0.8 AC=1
V_X100Y110VDD_X100Y110VSS X100Y110VDDDM X100Y110VSS 0
I_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VDDDM 0.8 AC=1
V_X110Y120VDD_X110Y120VSS X110Y120VDDDM X110Y120VSS 0
I_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VDDDM 0.8 AC=1
V_X110Y10VDD_X110Y10VSS X110Y10VDDDM X110Y10VSS 0
I_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VDDDM 0.8 AC=1
V_X110Y20VDD_X110Y20VSS X110Y20VDDDM X110Y20VSS 0
I_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VDDDM 0.8 AC=1
V_X110Y30VDD_X110Y30VSS X110Y30VDDDM X110Y30VSS 0
I_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VDDDM 0.8 AC=1
V_X110Y40VDD_X110Y40VSS X110Y40VDDDM X110Y40VSS 0
I_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VDDDM 0.8 AC=1
V_X110Y50VDD_X110Y50VSS X110Y50VDDDM X110Y50VSS 0
I_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VDDDM 0.8 AC=1
V_X110Y60VDD_X110Y60VSS X110Y60VDDDM X110Y60VSS 0
I_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VDDDM 0.8 AC=1
V_X110Y70VDD_X110Y70VSS X110Y70VDDDM X110Y70VSS 0
I_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VDDDM 0.8 AC=1
V_X110Y80VDD_X110Y80VSS X110Y80VDDDM X110Y80VSS 0
I_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VDDDM 0.8 AC=1
V_X110Y90VDD_X110Y90VSS X110Y90VDDDM X110Y90VSS 0
I_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VDDDM 0.8 AC=1
V_X110Y100VDD_X110Y100VSS X110Y100VDDDM X110Y100VSS 0
I_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VDDDM 0.8 AC=1
V_X110Y110VDD_X110Y110VSS X110Y110VDDDM X110Y110VSS 0
Rs1_1 VDD 11_1 0.027Ohm
Cp1_1 11_1 VSS 131.33333333333331nF
Rs2_1 11_1 12_1 0.027Ohm
Cp2_1 12_1 VSS 213.33333333333331nF
Fs_1 12_1 VSS V_X60Y60VDD_X60Y60VSS 3.0
Rg_1 VSS X60Y60VSS 0.025Ohm
Es_1 13_1 X60Y60VSS VDD VSS 0.3333333333333333
Rs3_1 13_1 14_1 0.009Ohm
Cp3_1 14_1 X60Y60VSS 394nF
Rs4_1 14_1 X60Y60VDD 0.009Ohm
Cp4_1 X60Y60VDD X60Y60VSS 640nF
.ends dut
XRegulator0 VDD0 VSS0 Regulator
Rgnd VSS0 0 0
XPcbModelLumped0 VDD0 VSS0 VDD1 VSS1 PcbModelLumped
XChipPackage1 VDD1 VSS1 VDD2 VSS2 ChipPackage
XChipBump2 VDD2 VSS2 VDD3 VSS3 ChipBump
Xdut3 VDD3 VSS3 dut


# case 1 feedback
.title 20200622-105330
.option rshunt = 1.0e12
.subckt PcbBuckConverter VDD VSS
C1 VDD 12 2340uF
R1 12 13 0Ohm
L1 13 VSS 0nH
C2 VDD 22 0uF
R2 22 23 1000000000000.0Ohm
L2 23 VSS 0nH
Ls VDD 31 0.33uH
Rs 31 32 20mOhm
Vs 32 VSS 1.1
.ends PcbBuckConverter

.subckt PcbModelLumped VDD1 VSS1 VDD2 VSS2
Rs1 VDD1 11 1000mOhm
Ls1 11 VDD2 0nH
Rs2 VSS1 21 1000mOhm
Ls2 21 VSS2 0nH
Rp VDD2 VDD2M 0mOhm
Cp VDD2M VSS2 0uF
.ends PcbModelLumped

.subckt dut VDD VSS
R_X10Y10VDD_X20Y10VDD X10Y10VDD X15Y10VDD 25mOhm
L_X10Y10VDD_X20Y10VDD X15Y10VDD X20Y10VDD 2.91e-06nH
R_X10Y10VSS_X20Y10VSS X10Y10VSS X15Y10VSS 25mOhm
L_X10Y10VSS_X20Y10VSS X15Y10VSS X20Y10VSS 2.91e-06nH
R_X20Y10VDD_X30Y10VDD X20Y10VDD X25Y10VDD 25mOhm
L_X20Y10VDD_X30Y10VDD X25Y10VDD X30Y10VDD 2.91e-06nH
R_X20Y10VSS_X30Y10VSS X20Y10VSS X25Y10VSS 25mOhm
L_X20Y10VSS_X30Y10VSS X25Y10VSS X30Y10VSS 2.91e-06nH
R_X30Y10VDD_X40Y10VDD X30Y10VDD X35Y10VDD 25mOhm
L_X30Y10VDD_X40Y10VDD X35Y10VDD X40Y10VDD 2.91e-06nH
R_X30Y10VSS_X40Y10VSS X30Y10VSS X35Y10VSS 25mOhm
L_X30Y10VSS_X40Y10VSS X35Y10VSS X40Y10VSS 2.91e-06nH
R_X40Y10VDD_X50Y10VDD X40Y10VDD X45Y10VDD 25mOhm
L_X40Y10VDD_X50Y10VDD X45Y10VDD X50Y10VDD 2.91e-06nH
R_X40Y10VSS_X50Y10VSS X40Y10VSS X45Y10VSS 25mOhm
L_X40Y10VSS_X50Y10VSS X45Y10VSS X50Y10VSS 2.91e-06nH
R_X50Y10VDD_X60Y10VDD X50Y10VDD X55Y10VDD 25mOhm
L_X50Y10VDD_X60Y10VDD X55Y10VDD X60Y10VDD 2.91e-06nH
R_X50Y10VSS_X60Y10VSS X50Y10VSS X55Y10VSS 25mOhm
L_X50Y10VSS_X60Y10VSS X55Y10VSS X60Y10VSS 2.91e-06nH
R_X60Y10VDD_X70Y10VDD X60Y10VDD X65Y10VDD 25mOhm
L_X60Y10VDD_X70Y10VDD X65Y10VDD X70Y10VDD 2.91e-06nH
R_X60Y10VSS_X70Y10VSS X60Y10VSS X65Y10VSS 25mOhm
L_X60Y10VSS_X70Y10VSS X65Y10VSS X70Y10VSS 2.91e-06nH
R_X70Y10VDD_X80Y10VDD X70Y10VDD X75Y10VDD 25mOhm
L_X70Y10VDD_X80Y10VDD X75Y10VDD X80Y10VDD 2.91e-06nH
R_X70Y10VSS_X80Y10VSS X70Y10VSS X75Y10VSS 25mOhm
L_X70Y10VSS_X80Y10VSS X75Y10VSS X80Y10VSS 2.91e-06nH
R_X80Y10VDD_X90Y10VDD X80Y10VDD X85Y10VDD 25mOhm
L_X80Y10VDD_X90Y10VDD X85Y10VDD X90Y10VDD 2.91e-06nH
R_X80Y10VSS_X90Y10VSS X80Y10VSS X85Y10VSS 25mOhm
L_X80Y10VSS_X90Y10VSS X85Y10VSS X90Y10VSS 2.91e-06nH
R_X90Y10VDD_X100Y10VDD X90Y10VDD X95Y10VDD 25mOhm
L_X90Y10VDD_X100Y10VDD X95Y10VDD X100Y10VDD 2.91e-06nH
R_X90Y10VSS_X100Y10VSS X90Y10VSS X95Y10VSS 25mOhm
L_X90Y10VSS_X100Y10VSS X95Y10VSS X100Y10VSS 2.91e-06nH
R_X100Y10VDD_X110Y10VDD X100Y10VDD X105Y10VDD 25mOhm
L_X100Y10VDD_X110Y10VDD X105Y10VDD X110Y10VDD 2.91e-06nH
R_X100Y10VSS_X110Y10VSS X100Y10VSS X105Y10VSS 25mOhm
L_X100Y10VSS_X110Y10VSS X105Y10VSS X110Y10VSS 2.91e-06nH
R_X110Y10VDD_X120Y10VDD X110Y10VDD X115Y10VDD 25mOhm
L_X110Y10VDD_X120Y10VDD X115Y10VDD X120Y10VDD 2.91e-06nH
R_X110Y10VSS_X120Y10VSS X110Y10VSS X115Y10VSS 25mOhm
L_X110Y10VSS_X120Y10VSS X115Y10VSS X120Y10VSS 2.91e-06nH
R_X10Y20VDD_X20Y20VDD X10Y20VDD X15Y20VDD 25mOhm
L_X10Y20VDD_X20Y20VDD X15Y20VDD X20Y20VDD 2.91e-06nH
R_X10Y20VSS_X20Y20VSS X10Y20VSS X15Y20VSS 25mOhm
L_X10Y20VSS_X20Y20VSS X15Y20VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X30Y20VDD X20Y20VDD X25Y20VDD 25mOhm
L_X20Y20VDD_X30Y20VDD X25Y20VDD X30Y20VDD 2.91e-06nH
R_X20Y20VSS_X30Y20VSS X20Y20VSS X25Y20VSS 25mOhm
L_X20Y20VSS_X30Y20VSS X25Y20VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X40Y20VDD X30Y20VDD X35Y20VDD 25mOhm
L_X30Y20VDD_X40Y20VDD X35Y20VDD X40Y20VDD 2.91e-06nH
R_X30Y20VSS_X40Y20VSS X30Y20VSS X35Y20VSS 25mOhm
L_X30Y20VSS_X40Y20VSS X35Y20VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X50Y20VDD X40Y20VDD X45Y20VDD 25mOhm
L_X40Y20VDD_X50Y20VDD X45Y20VDD X50Y20VDD 2.91e-06nH
R_X40Y20VSS_X50Y20VSS X40Y20VSS X45Y20VSS 25mOhm
L_X40Y20VSS_X50Y20VSS X45Y20VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X60Y20VDD X50Y20VDD X55Y20VDD 25mOhm
L_X50Y20VDD_X60Y20VDD X55Y20VDD X60Y20VDD 2.91e-06nH
R_X50Y20VSS_X60Y20VSS X50Y20VSS X55Y20VSS 25mOhm
L_X50Y20VSS_X60Y20VSS X55Y20VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X70Y20VDD X60Y20VDD X65Y20VDD 25mOhm
L_X60Y20VDD_X70Y20VDD X65Y20VDD X70Y20VDD 2.91e-06nH
R_X60Y20VSS_X70Y20VSS X60Y20VSS X65Y20VSS 25mOhm
L_X60Y20VSS_X70Y20VSS X65Y20VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X80Y20VDD X70Y20VDD X75Y20VDD 25mOhm
L_X70Y20VDD_X80Y20VDD X75Y20VDD X80Y20VDD 2.91e-06nH
R_X70Y20VSS_X80Y20VSS X70Y20VSS X75Y20VSS 25mOhm
L_X70Y20VSS_X80Y20VSS X75Y20VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X90Y20VDD X80Y20VDD X85Y20VDD 25mOhm
L_X80Y20VDD_X90Y20VDD X85Y20VDD X90Y20VDD 2.91e-06nH
R_X80Y20VSS_X90Y20VSS X80Y20VSS X85Y20VSS 25mOhm
L_X80Y20VSS_X90Y20VSS X85Y20VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X100Y20VDD X90Y20VDD X95Y20VDD 25mOhm
L_X90Y20VDD_X100Y20VDD X95Y20VDD X100Y20VDD 2.91e-06nH
R_X90Y20VSS_X100Y20VSS X90Y20VSS X95Y20VSS 25mOhm
L_X90Y20VSS_X100Y20VSS X95Y20VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X110Y20VDD X100Y20VDD X105Y20VDD 25mOhm
L_X100Y20VDD_X110Y20VDD X105Y20VDD X110Y20VDD 2.91e-06nH
R_X100Y20VSS_X110Y20VSS X100Y20VSS X105Y20VSS 25mOhm
L_X100Y20VSS_X110Y20VSS X105Y20VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X120Y20VDD X110Y20VDD X115Y20VDD 25mOhm
L_X110Y20VDD_X120Y20VDD X115Y20VDD X120Y20VDD 2.91e-06nH
R_X110Y20VSS_X120Y20VSS X110Y20VSS X115Y20VSS 25mOhm
L_X110Y20VSS_X120Y20VSS X115Y20VSS X120Y20VSS 2.91e-06nH
R_X10Y30VDD_X20Y30VDD X10Y30VDD X15Y30VDD 25mOhm
L_X10Y30VDD_X20Y30VDD X15Y30VDD X20Y30VDD 2.91e-06nH
R_X10Y30VSS_X20Y30VSS X10Y30VSS X15Y30VSS 25mOhm
L_X10Y30VSS_X20Y30VSS X15Y30VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X30Y30VDD X20Y30VDD X25Y30VDD 25mOhm
L_X20Y30VDD_X30Y30VDD X25Y30VDD X30Y30VDD 2.91e-06nH
R_X20Y30VSS_X30Y30VSS X20Y30VSS X25Y30VSS 25mOhm
L_X20Y30VSS_X30Y30VSS X25Y30VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X40Y30VDD X30Y30VDD X35Y30VDD 25mOhm
L_X30Y30VDD_X40Y30VDD X35Y30VDD X40Y30VDD 2.91e-06nH
R_X30Y30VSS_X40Y30VSS X30Y30VSS X35Y30VSS 25mOhm
L_X30Y30VSS_X40Y30VSS X35Y30VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X50Y30VDD X40Y30VDD X45Y30VDD 25mOhm
L_X40Y30VDD_X50Y30VDD X45Y30VDD X50Y30VDD 2.91e-06nH
R_X40Y30VSS_X50Y30VSS X40Y30VSS X45Y30VSS 25mOhm
L_X40Y30VSS_X50Y30VSS X45Y30VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X60Y30VDD X50Y30VDD X55Y30VDD 25mOhm
L_X50Y30VDD_X60Y30VDD X55Y30VDD X60Y30VDD 2.91e-06nH
R_X50Y30VSS_X60Y30VSS X50Y30VSS X55Y30VSS 25mOhm
L_X50Y30VSS_X60Y30VSS X55Y30VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X70Y30VDD X60Y30VDD X65Y30VDD 25mOhm
L_X60Y30VDD_X70Y30VDD X65Y30VDD X70Y30VDD 2.91e-06nH
R_X60Y30VSS_X70Y30VSS X60Y30VSS X65Y30VSS 25mOhm
L_X60Y30VSS_X70Y30VSS X65Y30VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X80Y30VDD X70Y30VDD X75Y30VDD 25mOhm
L_X70Y30VDD_X80Y30VDD X75Y30VDD X80Y30VDD 2.91e-06nH
R_X70Y30VSS_X80Y30VSS X70Y30VSS X75Y30VSS 25mOhm
L_X70Y30VSS_X80Y30VSS X75Y30VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X90Y30VDD X80Y30VDD X85Y30VDD 25mOhm
L_X80Y30VDD_X90Y30VDD X85Y30VDD X90Y30VDD 2.91e-06nH
R_X80Y30VSS_X90Y30VSS X80Y30VSS X85Y30VSS 25mOhm
L_X80Y30VSS_X90Y30VSS X85Y30VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X100Y30VDD X90Y30VDD X95Y30VDD 25mOhm
L_X90Y30VDD_X100Y30VDD X95Y30VDD X100Y30VDD 2.91e-06nH
R_X90Y30VSS_X100Y30VSS X90Y30VSS X95Y30VSS 25mOhm
L_X90Y30VSS_X100Y30VSS X95Y30VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X110Y30VDD X100Y30VDD X105Y30VDD 25mOhm
L_X100Y30VDD_X110Y30VDD X105Y30VDD X110Y30VDD 2.91e-06nH
R_X100Y30VSS_X110Y30VSS X100Y30VSS X105Y30VSS 25mOhm
L_X100Y30VSS_X110Y30VSS X105Y30VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X120Y30VDD X110Y30VDD X115Y30VDD 25mOhm
L_X110Y30VDD_X120Y30VDD X115Y30VDD X120Y30VDD 2.91e-06nH
R_X110Y30VSS_X120Y30VSS X110Y30VSS X115Y30VSS 25mOhm
L_X110Y30VSS_X120Y30VSS X115Y30VSS X120Y30VSS 2.91e-06nH
R_X10Y40VDD_X20Y40VDD X10Y40VDD X15Y40VDD 25mOhm
L_X10Y40VDD_X20Y40VDD X15Y40VDD X20Y40VDD 2.91e-06nH
R_X10Y40VSS_X20Y40VSS X10Y40VSS X15Y40VSS 25mOhm
L_X10Y40VSS_X20Y40VSS X15Y40VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X30Y40VDD X20Y40VDD X25Y40VDD 25mOhm
L_X20Y40VDD_X30Y40VDD X25Y40VDD X30Y40VDD 2.91e-06nH
R_X20Y40VSS_X30Y40VSS X20Y40VSS X25Y40VSS 25mOhm
L_X20Y40VSS_X30Y40VSS X25Y40VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X40Y40VDD X30Y40VDD X35Y40VDD 25mOhm
L_X30Y40VDD_X40Y40VDD X35Y40VDD X40Y40VDD 2.91e-06nH
R_X30Y40VSS_X40Y40VSS X30Y40VSS X35Y40VSS 25mOhm
L_X30Y40VSS_X40Y40VSS X35Y40VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X50Y40VDD X40Y40VDD X45Y40VDD 25mOhm
L_X40Y40VDD_X50Y40VDD X45Y40VDD X50Y40VDD 2.91e-06nH
R_X40Y40VSS_X50Y40VSS X40Y40VSS X45Y40VSS 25mOhm
L_X40Y40VSS_X50Y40VSS X45Y40VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X60Y40VDD X50Y40VDD X55Y40VDD 25mOhm
L_X50Y40VDD_X60Y40VDD X55Y40VDD X60Y40VDD 2.91e-06nH
R_X50Y40VSS_X60Y40VSS X50Y40VSS X55Y40VSS 25mOhm
L_X50Y40VSS_X60Y40VSS X55Y40VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X70Y40VDD X60Y40VDD X65Y40VDD 25mOhm
L_X60Y40VDD_X70Y40VDD X65Y40VDD X70Y40VDD 2.91e-06nH
R_X60Y40VSS_X70Y40VSS X60Y40VSS X65Y40VSS 25mOhm
L_X60Y40VSS_X70Y40VSS X65Y40VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X80Y40VDD X70Y40VDD X75Y40VDD 25mOhm
L_X70Y40VDD_X80Y40VDD X75Y40VDD X80Y40VDD 2.91e-06nH
R_X70Y40VSS_X80Y40VSS X70Y40VSS X75Y40VSS 25mOhm
L_X70Y40VSS_X80Y40VSS X75Y40VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X90Y40VDD X80Y40VDD X85Y40VDD 25mOhm
L_X80Y40VDD_X90Y40VDD X85Y40VDD X90Y40VDD 2.91e-06nH
R_X80Y40VSS_X90Y40VSS X80Y40VSS X85Y40VSS 25mOhm
L_X80Y40VSS_X90Y40VSS X85Y40VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X100Y40VDD X90Y40VDD X95Y40VDD 25mOhm
L_X90Y40VDD_X100Y40VDD X95Y40VDD X100Y40VDD 2.91e-06nH
R_X90Y40VSS_X100Y40VSS X90Y40VSS X95Y40VSS 25mOhm
L_X90Y40VSS_X100Y40VSS X95Y40VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X110Y40VDD X100Y40VDD X105Y40VDD 25mOhm
L_X100Y40VDD_X110Y40VDD X105Y40VDD X110Y40VDD 2.91e-06nH
R_X100Y40VSS_X110Y40VSS X100Y40VSS X105Y40VSS 25mOhm
L_X100Y40VSS_X110Y40VSS X105Y40VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X120Y40VDD X110Y40VDD X115Y40VDD 25mOhm
L_X110Y40VDD_X120Y40VDD X115Y40VDD X120Y40VDD 2.91e-06nH
R_X110Y40VSS_X120Y40VSS X110Y40VSS X115Y40VSS 25mOhm
L_X110Y40VSS_X120Y40VSS X115Y40VSS X120Y40VSS 2.91e-06nH
R_X10Y50VDD_X20Y50VDD X10Y50VDD X15Y50VDD 25mOhm
L_X10Y50VDD_X20Y50VDD X15Y50VDD X20Y50VDD 2.91e-06nH
R_X10Y50VSS_X20Y50VSS X10Y50VSS X15Y50VSS 25mOhm
L_X10Y50VSS_X20Y50VSS X15Y50VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X30Y50VDD X20Y50VDD X25Y50VDD 25mOhm
L_X20Y50VDD_X30Y50VDD X25Y50VDD X30Y50VDD 2.91e-06nH
R_X20Y50VSS_X30Y50VSS X20Y50VSS X25Y50VSS 25mOhm
L_X20Y50VSS_X30Y50VSS X25Y50VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X40Y50VDD X30Y50VDD X35Y50VDD 25mOhm
L_X30Y50VDD_X40Y50VDD X35Y50VDD X40Y50VDD 2.91e-06nH
R_X30Y50VSS_X40Y50VSS X30Y50VSS X35Y50VSS 25mOhm
L_X30Y50VSS_X40Y50VSS X35Y50VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X50Y50VDD X40Y50VDD X45Y50VDD 25mOhm
L_X40Y50VDD_X50Y50VDD X45Y50VDD X50Y50VDD 2.91e-06nH
R_X40Y50VSS_X50Y50VSS X40Y50VSS X45Y50VSS 25mOhm
L_X40Y50VSS_X50Y50VSS X45Y50VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X60Y50VDD X50Y50VDD X55Y50VDD 25mOhm
L_X50Y50VDD_X60Y50VDD X55Y50VDD X60Y50VDD 2.91e-06nH
R_X50Y50VSS_X60Y50VSS X50Y50VSS X55Y50VSS 25mOhm
L_X50Y50VSS_X60Y50VSS X55Y50VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X70Y50VDD X60Y50VDD X65Y50VDD 25mOhm
L_X60Y50VDD_X70Y50VDD X65Y50VDD X70Y50VDD 2.91e-06nH
R_X60Y50VSS_X70Y50VSS X60Y50VSS X65Y50VSS 25mOhm
L_X60Y50VSS_X70Y50VSS X65Y50VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X80Y50VDD X70Y50VDD X75Y50VDD 25mOhm
L_X70Y50VDD_X80Y50VDD X75Y50VDD X80Y50VDD 2.91e-06nH
R_X70Y50VSS_X80Y50VSS X70Y50VSS X75Y50VSS 25mOhm
L_X70Y50VSS_X80Y50VSS X75Y50VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X90Y50VDD X80Y50VDD X85Y50VDD 25mOhm
L_X80Y50VDD_X90Y50VDD X85Y50VDD X90Y50VDD 2.91e-06nH
R_X80Y50VSS_X90Y50VSS X80Y50VSS X85Y50VSS 25mOhm
L_X80Y50VSS_X90Y50VSS X85Y50VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X100Y50VDD X90Y50VDD X95Y50VDD 25mOhm
L_X90Y50VDD_X100Y50VDD X95Y50VDD X100Y50VDD 2.91e-06nH
R_X90Y50VSS_X100Y50VSS X90Y50VSS X95Y50VSS 25mOhm
L_X90Y50VSS_X100Y50VSS X95Y50VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X110Y50VDD X100Y50VDD X105Y50VDD 25mOhm
L_X100Y50VDD_X110Y50VDD X105Y50VDD X110Y50VDD 2.91e-06nH
R_X100Y50VSS_X110Y50VSS X100Y50VSS X105Y50VSS 25mOhm
L_X100Y50VSS_X110Y50VSS X105Y50VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X120Y50VDD X110Y50VDD X115Y50VDD 25mOhm
L_X110Y50VDD_X120Y50VDD X115Y50VDD X120Y50VDD 2.91e-06nH
R_X110Y50VSS_X120Y50VSS X110Y50VSS X115Y50VSS 25mOhm
L_X110Y50VSS_X120Y50VSS X115Y50VSS X120Y50VSS 2.91e-06nH
R_X10Y60VDD_X20Y60VDD X10Y60VDD X15Y60VDD 25mOhm
L_X10Y60VDD_X20Y60VDD X15Y60VDD X20Y60VDD 2.91e-06nH
R_X10Y60VSS_X20Y60VSS X10Y60VSS X15Y60VSS 25mOhm
L_X10Y60VSS_X20Y60VSS X15Y60VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X30Y60VDD X20Y60VDD X25Y60VDD 25mOhm
L_X20Y60VDD_X30Y60VDD X25Y60VDD X30Y60VDD 2.91e-06nH
R_X20Y60VSS_X30Y60VSS X20Y60VSS X25Y60VSS 25mOhm
L_X20Y60VSS_X30Y60VSS X25Y60VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X40Y60VDD X30Y60VDD X35Y60VDD 25mOhm
L_X30Y60VDD_X40Y60VDD X35Y60VDD X40Y60VDD 2.91e-06nH
R_X30Y60VSS_X40Y60VSS X30Y60VSS X35Y60VSS 25mOhm
L_X30Y60VSS_X40Y60VSS X35Y60VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X50Y60VDD X40Y60VDD X45Y60VDD 25mOhm
L_X40Y60VDD_X50Y60VDD X45Y60VDD X50Y60VDD 2.91e-06nH
R_X40Y60VSS_X50Y60VSS X40Y60VSS X45Y60VSS 25mOhm
L_X40Y60VSS_X50Y60VSS X45Y60VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X60Y60VDD X50Y60VDD X55Y60VDD 25mOhm
L_X50Y60VDD_X60Y60VDD X55Y60VDD X60Y60VDD 2.91e-06nH
R_X50Y60VSS_X60Y60VSS X50Y60VSS X55Y60VSS 25mOhm
L_X50Y60VSS_X60Y60VSS X55Y60VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X70Y60VDD X60Y60VDD X65Y60VDD 25mOhm
L_X60Y60VDD_X70Y60VDD X65Y60VDD X70Y60VDD 2.91e-06nH
R_X60Y60VSS_X70Y60VSS X60Y60VSS X65Y60VSS 25mOhm
L_X60Y60VSS_X70Y60VSS X65Y60VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X80Y60VDD X70Y60VDD X75Y60VDD 25mOhm
L_X70Y60VDD_X80Y60VDD X75Y60VDD X80Y60VDD 2.91e-06nH
R_X70Y60VSS_X80Y60VSS X70Y60VSS X75Y60VSS 25mOhm
L_X70Y60VSS_X80Y60VSS X75Y60VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X90Y60VDD X80Y60VDD X85Y60VDD 25mOhm
L_X80Y60VDD_X90Y60VDD X85Y60VDD X90Y60VDD 2.91e-06nH
R_X80Y60VSS_X90Y60VSS X80Y60VSS X85Y60VSS 25mOhm
L_X80Y60VSS_X90Y60VSS X85Y60VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X100Y60VDD X90Y60VDD X95Y60VDD 25mOhm
L_X90Y60VDD_X100Y60VDD X95Y60VDD X100Y60VDD 2.91e-06nH
R_X90Y60VSS_X100Y60VSS X90Y60VSS X95Y60VSS 25mOhm
L_X90Y60VSS_X100Y60VSS X95Y60VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X110Y60VDD X100Y60VDD X105Y60VDD 25mOhm
L_X100Y60VDD_X110Y60VDD X105Y60VDD X110Y60VDD 2.91e-06nH
R_X100Y60VSS_X110Y60VSS X100Y60VSS X105Y60VSS 25mOhm
L_X100Y60VSS_X110Y60VSS X105Y60VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X120Y60VDD X110Y60VDD X115Y60VDD 25mOhm
L_X110Y60VDD_X120Y60VDD X115Y60VDD X120Y60VDD 2.91e-06nH
R_X110Y60VSS_X120Y60VSS X110Y60VSS X115Y60VSS 25mOhm
L_X110Y60VSS_X120Y60VSS X115Y60VSS X120Y60VSS 2.91e-06nH
R_X10Y70VDD_X20Y70VDD X10Y70VDD X15Y70VDD 25mOhm
L_X10Y70VDD_X20Y70VDD X15Y70VDD X20Y70VDD 2.91e-06nH
R_X10Y70VSS_X20Y70VSS X10Y70VSS X15Y70VSS 25mOhm
L_X10Y70VSS_X20Y70VSS X15Y70VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X30Y70VDD X20Y70VDD X25Y70VDD 25mOhm
L_X20Y70VDD_X30Y70VDD X25Y70VDD X30Y70VDD 2.91e-06nH
R_X20Y70VSS_X30Y70VSS X20Y70VSS X25Y70VSS 25mOhm
L_X20Y70VSS_X30Y70VSS X25Y70VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X40Y70VDD X30Y70VDD X35Y70VDD 25mOhm
L_X30Y70VDD_X40Y70VDD X35Y70VDD X40Y70VDD 2.91e-06nH
R_X30Y70VSS_X40Y70VSS X30Y70VSS X35Y70VSS 25mOhm
L_X30Y70VSS_X40Y70VSS X35Y70VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X50Y70VDD X40Y70VDD X45Y70VDD 25mOhm
L_X40Y70VDD_X50Y70VDD X45Y70VDD X50Y70VDD 2.91e-06nH
R_X40Y70VSS_X50Y70VSS X40Y70VSS X45Y70VSS 25mOhm
L_X40Y70VSS_X50Y70VSS X45Y70VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X60Y70VDD X50Y70VDD X55Y70VDD 25mOhm
L_X50Y70VDD_X60Y70VDD X55Y70VDD X60Y70VDD 2.91e-06nH
R_X50Y70VSS_X60Y70VSS X50Y70VSS X55Y70VSS 25mOhm
L_X50Y70VSS_X60Y70VSS X55Y70VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X70Y70VDD X60Y70VDD X65Y70VDD 25mOhm
L_X60Y70VDD_X70Y70VDD X65Y70VDD X70Y70VDD 2.91e-06nH
R_X60Y70VSS_X70Y70VSS X60Y70VSS X65Y70VSS 25mOhm
L_X60Y70VSS_X70Y70VSS X65Y70VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X80Y70VDD X70Y70VDD X75Y70VDD 25mOhm
L_X70Y70VDD_X80Y70VDD X75Y70VDD X80Y70VDD 2.91e-06nH
R_X70Y70VSS_X80Y70VSS X70Y70VSS X75Y70VSS 25mOhm
L_X70Y70VSS_X80Y70VSS X75Y70VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X90Y70VDD X80Y70VDD X85Y70VDD 25mOhm
L_X80Y70VDD_X90Y70VDD X85Y70VDD X90Y70VDD 2.91e-06nH
R_X80Y70VSS_X90Y70VSS X80Y70VSS X85Y70VSS 25mOhm
L_X80Y70VSS_X90Y70VSS X85Y70VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X100Y70VDD X90Y70VDD X95Y70VDD 25mOhm
L_X90Y70VDD_X100Y70VDD X95Y70VDD X100Y70VDD 2.91e-06nH
R_X90Y70VSS_X100Y70VSS X90Y70VSS X95Y70VSS 25mOhm
L_X90Y70VSS_X100Y70VSS X95Y70VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X110Y70VDD X100Y70VDD X105Y70VDD 25mOhm
L_X100Y70VDD_X110Y70VDD X105Y70VDD X110Y70VDD 2.91e-06nH
R_X100Y70VSS_X110Y70VSS X100Y70VSS X105Y70VSS 25mOhm
L_X100Y70VSS_X110Y70VSS X105Y70VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X120Y70VDD X110Y70VDD X115Y70VDD 25mOhm
L_X110Y70VDD_X120Y70VDD X115Y70VDD X120Y70VDD 2.91e-06nH
R_X110Y70VSS_X120Y70VSS X110Y70VSS X115Y70VSS 25mOhm
L_X110Y70VSS_X120Y70VSS X115Y70VSS X120Y70VSS 2.91e-06nH
R_X10Y80VDD_X20Y80VDD X10Y80VDD X15Y80VDD 25mOhm
L_X10Y80VDD_X20Y80VDD X15Y80VDD X20Y80VDD 2.91e-06nH
R_X10Y80VSS_X20Y80VSS X10Y80VSS X15Y80VSS 25mOhm
L_X10Y80VSS_X20Y80VSS X15Y80VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X30Y80VDD X20Y80VDD X25Y80VDD 25mOhm
L_X20Y80VDD_X30Y80VDD X25Y80VDD X30Y80VDD 2.91e-06nH
R_X20Y80VSS_X30Y80VSS X20Y80VSS X25Y80VSS 25mOhm
L_X20Y80VSS_X30Y80VSS X25Y80VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X40Y80VDD X30Y80VDD X35Y80VDD 25mOhm
L_X30Y80VDD_X40Y80VDD X35Y80VDD X40Y80VDD 2.91e-06nH
R_X30Y80VSS_X40Y80VSS X30Y80VSS X35Y80VSS 25mOhm
L_X30Y80VSS_X40Y80VSS X35Y80VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X50Y80VDD X40Y80VDD X45Y80VDD 25mOhm
L_X40Y80VDD_X50Y80VDD X45Y80VDD X50Y80VDD 2.91e-06nH
R_X40Y80VSS_X50Y80VSS X40Y80VSS X45Y80VSS 25mOhm
L_X40Y80VSS_X50Y80VSS X45Y80VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X60Y80VDD X50Y80VDD X55Y80VDD 25mOhm
L_X50Y80VDD_X60Y80VDD X55Y80VDD X60Y80VDD 2.91e-06nH
R_X50Y80VSS_X60Y80VSS X50Y80VSS X55Y80VSS 25mOhm
L_X50Y80VSS_X60Y80VSS X55Y80VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X70Y80VDD X60Y80VDD X65Y80VDD 25mOhm
L_X60Y80VDD_X70Y80VDD X65Y80VDD X70Y80VDD 2.91e-06nH
R_X60Y80VSS_X70Y80VSS X60Y80VSS X65Y80VSS 25mOhm
L_X60Y80VSS_X70Y80VSS X65Y80VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X80Y80VDD X70Y80VDD X75Y80VDD 25mOhm
L_X70Y80VDD_X80Y80VDD X75Y80VDD X80Y80VDD 2.91e-06nH
R_X70Y80VSS_X80Y80VSS X70Y80VSS X75Y80VSS 25mOhm
L_X70Y80VSS_X80Y80VSS X75Y80VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X90Y80VDD X80Y80VDD X85Y80VDD 25mOhm
L_X80Y80VDD_X90Y80VDD X85Y80VDD X90Y80VDD 2.91e-06nH
R_X80Y80VSS_X90Y80VSS X80Y80VSS X85Y80VSS 25mOhm
L_X80Y80VSS_X90Y80VSS X85Y80VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X100Y80VDD X90Y80VDD X95Y80VDD 25mOhm
L_X90Y80VDD_X100Y80VDD X95Y80VDD X100Y80VDD 2.91e-06nH
R_X90Y80VSS_X100Y80VSS X90Y80VSS X95Y80VSS 25mOhm
L_X90Y80VSS_X100Y80VSS X95Y80VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X110Y80VDD X100Y80VDD X105Y80VDD 25mOhm
L_X100Y80VDD_X110Y80VDD X105Y80VDD X110Y80VDD 2.91e-06nH
R_X100Y80VSS_X110Y80VSS X100Y80VSS X105Y80VSS 25mOhm
L_X100Y80VSS_X110Y80VSS X105Y80VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X120Y80VDD X110Y80VDD X115Y80VDD 25mOhm
L_X110Y80VDD_X120Y80VDD X115Y80VDD X120Y80VDD 2.91e-06nH
R_X110Y80VSS_X120Y80VSS X110Y80VSS X115Y80VSS 25mOhm
L_X110Y80VSS_X120Y80VSS X115Y80VSS X120Y80VSS 2.91e-06nH
R_X10Y90VDD_X20Y90VDD X10Y90VDD X15Y90VDD 25mOhm
L_X10Y90VDD_X20Y90VDD X15Y90VDD X20Y90VDD 2.91e-06nH
R_X10Y90VSS_X20Y90VSS X10Y90VSS X15Y90VSS 25mOhm
L_X10Y90VSS_X20Y90VSS X15Y90VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X30Y90VDD X20Y90VDD X25Y90VDD 25mOhm
L_X20Y90VDD_X30Y90VDD X25Y90VDD X30Y90VDD 2.91e-06nH
R_X20Y90VSS_X30Y90VSS X20Y90VSS X25Y90VSS 25mOhm
L_X20Y90VSS_X30Y90VSS X25Y90VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X40Y90VDD X30Y90VDD X35Y90VDD 25mOhm
L_X30Y90VDD_X40Y90VDD X35Y90VDD X40Y90VDD 2.91e-06nH
R_X30Y90VSS_X40Y90VSS X30Y90VSS X35Y90VSS 25mOhm
L_X30Y90VSS_X40Y90VSS X35Y90VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X50Y90VDD X40Y90VDD X45Y90VDD 25mOhm
L_X40Y90VDD_X50Y90VDD X45Y90VDD X50Y90VDD 2.91e-06nH
R_X40Y90VSS_X50Y90VSS X40Y90VSS X45Y90VSS 25mOhm
L_X40Y90VSS_X50Y90VSS X45Y90VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X60Y90VDD X50Y90VDD X55Y90VDD 25mOhm
L_X50Y90VDD_X60Y90VDD X55Y90VDD X60Y90VDD 2.91e-06nH
R_X50Y90VSS_X60Y90VSS X50Y90VSS X55Y90VSS 25mOhm
L_X50Y90VSS_X60Y90VSS X55Y90VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X70Y90VDD X60Y90VDD X65Y90VDD 25mOhm
L_X60Y90VDD_X70Y90VDD X65Y90VDD X70Y90VDD 2.91e-06nH
R_X60Y90VSS_X70Y90VSS X60Y90VSS X65Y90VSS 25mOhm
L_X60Y90VSS_X70Y90VSS X65Y90VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X80Y90VDD X70Y90VDD X75Y90VDD 25mOhm
L_X70Y90VDD_X80Y90VDD X75Y90VDD X80Y90VDD 2.91e-06nH
R_X70Y90VSS_X80Y90VSS X70Y90VSS X75Y90VSS 25mOhm
L_X70Y90VSS_X80Y90VSS X75Y90VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X90Y90VDD X80Y90VDD X85Y90VDD 25mOhm
L_X80Y90VDD_X90Y90VDD X85Y90VDD X90Y90VDD 2.91e-06nH
R_X80Y90VSS_X90Y90VSS X80Y90VSS X85Y90VSS 25mOhm
L_X80Y90VSS_X90Y90VSS X85Y90VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X100Y90VDD X90Y90VDD X95Y90VDD 25mOhm
L_X90Y90VDD_X100Y90VDD X95Y90VDD X100Y90VDD 2.91e-06nH
R_X90Y90VSS_X100Y90VSS X90Y90VSS X95Y90VSS 25mOhm
L_X90Y90VSS_X100Y90VSS X95Y90VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X110Y90VDD X100Y90VDD X105Y90VDD 25mOhm
L_X100Y90VDD_X110Y90VDD X105Y90VDD X110Y90VDD 2.91e-06nH
R_X100Y90VSS_X110Y90VSS X100Y90VSS X105Y90VSS 25mOhm
L_X100Y90VSS_X110Y90VSS X105Y90VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X120Y90VDD X110Y90VDD X115Y90VDD 25mOhm
L_X110Y90VDD_X120Y90VDD X115Y90VDD X120Y90VDD 2.91e-06nH
R_X110Y90VSS_X120Y90VSS X110Y90VSS X115Y90VSS 25mOhm
L_X110Y90VSS_X120Y90VSS X115Y90VSS X120Y90VSS 2.91e-06nH
R_X10Y100VDD_X20Y100VDD X10Y100VDD X15Y100VDD 25mOhm
L_X10Y100VDD_X20Y100VDD X15Y100VDD X20Y100VDD 2.91e-06nH
R_X10Y100VSS_X20Y100VSS X10Y100VSS X15Y100VSS 25mOhm
L_X10Y100VSS_X20Y100VSS X15Y100VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X30Y100VDD X20Y100VDD X25Y100VDD 25mOhm
L_X20Y100VDD_X30Y100VDD X25Y100VDD X30Y100VDD 2.91e-06nH
R_X20Y100VSS_X30Y100VSS X20Y100VSS X25Y100VSS 25mOhm
L_X20Y100VSS_X30Y100VSS X25Y100VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X40Y100VDD X30Y100VDD X35Y100VDD 25mOhm
L_X30Y100VDD_X40Y100VDD X35Y100VDD X40Y100VDD 2.91e-06nH
R_X30Y100VSS_X40Y100VSS X30Y100VSS X35Y100VSS 25mOhm
L_X30Y100VSS_X40Y100VSS X35Y100VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X50Y100VDD X40Y100VDD X45Y100VDD 25mOhm
L_X40Y100VDD_X50Y100VDD X45Y100VDD X50Y100VDD 2.91e-06nH
R_X40Y100VSS_X50Y100VSS X40Y100VSS X45Y100VSS 25mOhm
L_X40Y100VSS_X50Y100VSS X45Y100VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X60Y100VDD X50Y100VDD X55Y100VDD 25mOhm
L_X50Y100VDD_X60Y100VDD X55Y100VDD X60Y100VDD 2.91e-06nH
R_X50Y100VSS_X60Y100VSS X50Y100VSS X55Y100VSS 25mOhm
L_X50Y100VSS_X60Y100VSS X55Y100VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X70Y100VDD X60Y100VDD X65Y100VDD 25mOhm
L_X60Y100VDD_X70Y100VDD X65Y100VDD X70Y100VDD 2.91e-06nH
R_X60Y100VSS_X70Y100VSS X60Y100VSS X65Y100VSS 25mOhm
L_X60Y100VSS_X70Y100VSS X65Y100VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X80Y100VDD X70Y100VDD X75Y100VDD 25mOhm
L_X70Y100VDD_X80Y100VDD X75Y100VDD X80Y100VDD 2.91e-06nH
R_X70Y100VSS_X80Y100VSS X70Y100VSS X75Y100VSS 25mOhm
L_X70Y100VSS_X80Y100VSS X75Y100VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X90Y100VDD X80Y100VDD X85Y100VDD 25mOhm
L_X80Y100VDD_X90Y100VDD X85Y100VDD X90Y100VDD 2.91e-06nH
R_X80Y100VSS_X90Y100VSS X80Y100VSS X85Y100VSS 25mOhm
L_X80Y100VSS_X90Y100VSS X85Y100VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X100Y100VDD X90Y100VDD X95Y100VDD 25mOhm
L_X90Y100VDD_X100Y100VDD X95Y100VDD X100Y100VDD 2.91e-06nH
R_X90Y100VSS_X100Y100VSS X90Y100VSS X95Y100VSS 25mOhm
L_X90Y100VSS_X100Y100VSS X95Y100VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X110Y100VDD X100Y100VDD X105Y100VDD 25mOhm
L_X100Y100VDD_X110Y100VDD X105Y100VDD X110Y100VDD 2.91e-06nH
R_X100Y100VSS_X110Y100VSS X100Y100VSS X105Y100VSS 25mOhm
L_X100Y100VSS_X110Y100VSS X105Y100VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X120Y100VDD X110Y100VDD X115Y100VDD 25mOhm
L_X110Y100VDD_X120Y100VDD X115Y100VDD X120Y100VDD 2.91e-06nH
R_X110Y100VSS_X120Y100VSS X110Y100VSS X115Y100VSS 25mOhm
L_X110Y100VSS_X120Y100VSS X115Y100VSS X120Y100VSS 2.91e-06nH
R_X10Y110VDD_X20Y110VDD X10Y110VDD X15Y110VDD 25mOhm
L_X10Y110VDD_X20Y110VDD X15Y110VDD X20Y110VDD 2.91e-06nH
R_X10Y110VSS_X20Y110VSS X10Y110VSS X15Y110VSS 25mOhm
L_X10Y110VSS_X20Y110VSS X15Y110VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X30Y110VDD X20Y110VDD X25Y110VDD 25mOhm
L_X20Y110VDD_X30Y110VDD X25Y110VDD X30Y110VDD 2.91e-06nH
R_X20Y110VSS_X30Y110VSS X20Y110VSS X25Y110VSS 25mOhm
L_X20Y110VSS_X30Y110VSS X25Y110VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X40Y110VDD X30Y110VDD X35Y110VDD 25mOhm
L_X30Y110VDD_X40Y110VDD X35Y110VDD X40Y110VDD 2.91e-06nH
R_X30Y110VSS_X40Y110VSS X30Y110VSS X35Y110VSS 25mOhm
L_X30Y110VSS_X40Y110VSS X35Y110VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X50Y110VDD X40Y110VDD X45Y110VDD 25mOhm
L_X40Y110VDD_X50Y110VDD X45Y110VDD X50Y110VDD 2.91e-06nH
R_X40Y110VSS_X50Y110VSS X40Y110VSS X45Y110VSS 25mOhm
L_X40Y110VSS_X50Y110VSS X45Y110VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X60Y110VDD X50Y110VDD X55Y110VDD 25mOhm
L_X50Y110VDD_X60Y110VDD X55Y110VDD X60Y110VDD 2.91e-06nH
R_X50Y110VSS_X60Y110VSS X50Y110VSS X55Y110VSS 25mOhm
L_X50Y110VSS_X60Y110VSS X55Y110VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X70Y110VDD X60Y110VDD X65Y110VDD 25mOhm
L_X60Y110VDD_X70Y110VDD X65Y110VDD X70Y110VDD 2.91e-06nH
R_X60Y110VSS_X70Y110VSS X60Y110VSS X65Y110VSS 25mOhm
L_X60Y110VSS_X70Y110VSS X65Y110VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X80Y110VDD X70Y110VDD X75Y110VDD 25mOhm
L_X70Y110VDD_X80Y110VDD X75Y110VDD X80Y110VDD 2.91e-06nH
R_X70Y110VSS_X80Y110VSS X70Y110VSS X75Y110VSS 25mOhm
L_X70Y110VSS_X80Y110VSS X75Y110VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X90Y110VDD X80Y110VDD X85Y110VDD 25mOhm
L_X80Y110VDD_X90Y110VDD X85Y110VDD X90Y110VDD 2.91e-06nH
R_X80Y110VSS_X90Y110VSS X80Y110VSS X85Y110VSS 25mOhm
L_X80Y110VSS_X90Y110VSS X85Y110VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X100Y110VDD X90Y110VDD X95Y110VDD 25mOhm
L_X90Y110VDD_X100Y110VDD X95Y110VDD X100Y110VDD 2.91e-06nH
R_X90Y110VSS_X100Y110VSS X90Y110VSS X95Y110VSS 25mOhm
L_X90Y110VSS_X100Y110VSS X95Y110VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X110Y110VDD X100Y110VDD X105Y110VDD 25mOhm
L_X100Y110VDD_X110Y110VDD X105Y110VDD X110Y110VDD 2.91e-06nH
R_X100Y110VSS_X110Y110VSS X100Y110VSS X105Y110VSS 25mOhm
L_X100Y110VSS_X110Y110VSS X105Y110VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X120Y110VDD X110Y110VDD X115Y110VDD 25mOhm
L_X110Y110VDD_X120Y110VDD X115Y110VDD X120Y110VDD 2.91e-06nH
R_X110Y110VSS_X120Y110VSS X110Y110VSS X115Y110VSS 25mOhm
L_X110Y110VSS_X120Y110VSS X115Y110VSS X120Y110VSS 2.91e-06nH
R_X10Y120VDD_X20Y120VDD X10Y120VDD X15Y120VDD 25mOhm
L_X10Y120VDD_X20Y120VDD X15Y120VDD X20Y120VDD 2.91e-06nH
R_X10Y120VSS_X20Y120VSS X10Y120VSS X15Y120VSS 25mOhm
L_X10Y120VSS_X20Y120VSS X15Y120VSS X20Y120VSS 2.91e-06nH
R_X20Y120VDD_X30Y120VDD X20Y120VDD X25Y120VDD 25mOhm
L_X20Y120VDD_X30Y120VDD X25Y120VDD X30Y120VDD 2.91e-06nH
R_X20Y120VSS_X30Y120VSS X20Y120VSS X25Y120VSS 25mOhm
L_X20Y120VSS_X30Y120VSS X25Y120VSS X30Y120VSS 2.91e-06nH
R_X30Y120VDD_X40Y120VDD X30Y120VDD X35Y120VDD 25mOhm
L_X30Y120VDD_X40Y120VDD X35Y120VDD X40Y120VDD 2.91e-06nH
R_X30Y120VSS_X40Y120VSS X30Y120VSS X35Y120VSS 25mOhm
L_X30Y120VSS_X40Y120VSS X35Y120VSS X40Y120VSS 2.91e-06nH
R_X40Y120VDD_X50Y120VDD X40Y120VDD X45Y120VDD 25mOhm
L_X40Y120VDD_X50Y120VDD X45Y120VDD X50Y120VDD 2.91e-06nH
R_X40Y120VSS_X50Y120VSS X40Y120VSS X45Y120VSS 25mOhm
L_X40Y120VSS_X50Y120VSS X45Y120VSS X50Y120VSS 2.91e-06nH
R_X50Y120VDD_X60Y120VDD X50Y120VDD X55Y120VDD 25mOhm
L_X50Y120VDD_X60Y120VDD X55Y120VDD X60Y120VDD 2.91e-06nH
R_X50Y120VSS_X60Y120VSS X50Y120VSS X55Y120VSS 25mOhm
L_X50Y120VSS_X60Y120VSS X55Y120VSS X60Y120VSS 2.91e-06nH
R_X60Y120VDD_X70Y120VDD X60Y120VDD X65Y120VDD 25mOhm
L_X60Y120VDD_X70Y120VDD X65Y120VDD X70Y120VDD 2.91e-06nH
R_X60Y120VSS_X70Y120VSS X60Y120VSS X65Y120VSS 25mOhm
L_X60Y120VSS_X70Y120VSS X65Y120VSS X70Y120VSS 2.91e-06nH
R_X70Y120VDD_X80Y120VDD X70Y120VDD X75Y120VDD 25mOhm
L_X70Y120VDD_X80Y120VDD X75Y120VDD X80Y120VDD 2.91e-06nH
R_X70Y120VSS_X80Y120VSS X70Y120VSS X75Y120VSS 25mOhm
L_X70Y120VSS_X80Y120VSS X75Y120VSS X80Y120VSS 2.91e-06nH
R_X80Y120VDD_X90Y120VDD X80Y120VDD X85Y120VDD 25mOhm
L_X80Y120VDD_X90Y120VDD X85Y120VDD X90Y120VDD 2.91e-06nH
R_X80Y120VSS_X90Y120VSS X80Y120VSS X85Y120VSS 25mOhm
L_X80Y120VSS_X90Y120VSS X85Y120VSS X90Y120VSS 2.91e-06nH
R_X90Y120VDD_X100Y120VDD X90Y120VDD X95Y120VDD 25mOhm
L_X90Y120VDD_X100Y120VDD X95Y120VDD X100Y120VDD 2.91e-06nH
R_X90Y120VSS_X100Y120VSS X90Y120VSS X95Y120VSS 25mOhm
L_X90Y120VSS_X100Y120VSS X95Y120VSS X100Y120VSS 2.91e-06nH
R_X100Y120VDD_X110Y120VDD X100Y120VDD X105Y120VDD 25mOhm
L_X100Y120VDD_X110Y120VDD X105Y120VDD X110Y120VDD 2.91e-06nH
R_X100Y120VSS_X110Y120VSS X100Y120VSS X105Y120VSS 25mOhm
L_X100Y120VSS_X110Y120VSS X105Y120VSS X110Y120VSS 2.91e-06nH
R_X110Y120VDD_X120Y120VDD X110Y120VDD X115Y120VDD 25mOhm
L_X110Y120VDD_X120Y120VDD X115Y120VDD X120Y120VDD 2.91e-06nH
R_X110Y120VSS_X120Y120VSS X110Y120VSS X115Y120VSS 25mOhm
L_X110Y120VSS_X120Y120VSS X115Y120VSS X120Y120VSS 2.91e-06nH
R_X10Y10VDD_X10Y20VDD X10Y10VDD X10Y15VDD 25mOhm
L_X10Y10VDD_X10Y20VDD X10Y15VDD X10Y20VDD 2.91e-06nH
R_X10Y10VSS_X10Y20VSS X10Y10VSS X10Y15VSS 25mOhm
L_X10Y10VSS_X10Y20VSS X10Y15VSS X10Y20VSS 2.91e-06nH
R_X10Y20VDD_X10Y30VDD X10Y20VDD X10Y25VDD 25mOhm
L_X10Y20VDD_X10Y30VDD X10Y25VDD X10Y30VDD 2.91e-06nH
R_X10Y20VSS_X10Y30VSS X10Y20VSS X10Y25VSS 25mOhm
L_X10Y20VSS_X10Y30VSS X10Y25VSS X10Y30VSS 2.91e-06nH
R_X10Y30VDD_X10Y40VDD X10Y30VDD X10Y35VDD 25mOhm
L_X10Y30VDD_X10Y40VDD X10Y35VDD X10Y40VDD 2.91e-06nH
R_X10Y30VSS_X10Y40VSS X10Y30VSS X10Y35VSS 25mOhm
L_X10Y30VSS_X10Y40VSS X10Y35VSS X10Y40VSS 2.91e-06nH
R_X10Y40VDD_X10Y50VDD X10Y40VDD X10Y45VDD 25mOhm
L_X10Y40VDD_X10Y50VDD X10Y45VDD X10Y50VDD 2.91e-06nH
R_X10Y40VSS_X10Y50VSS X10Y40VSS X10Y45VSS 25mOhm
L_X10Y40VSS_X10Y50VSS X10Y45VSS X10Y50VSS 2.91e-06nH
R_X10Y50VDD_X10Y60VDD X10Y50VDD X10Y55VDD 25mOhm
L_X10Y50VDD_X10Y60VDD X10Y55VDD X10Y60VDD 2.91e-06nH
R_X10Y50VSS_X10Y60VSS X10Y50VSS X10Y55VSS 25mOhm
L_X10Y50VSS_X10Y60VSS X10Y55VSS X10Y60VSS 2.91e-06nH
R_X10Y60VDD_X10Y70VDD X10Y60VDD X10Y65VDD 25mOhm
L_X10Y60VDD_X10Y70VDD X10Y65VDD X10Y70VDD 2.91e-06nH
R_X10Y60VSS_X10Y70VSS X10Y60VSS X10Y65VSS 25mOhm
L_X10Y60VSS_X10Y70VSS X10Y65VSS X10Y70VSS 2.91e-06nH
R_X10Y70VDD_X10Y80VDD X10Y70VDD X10Y75VDD 25mOhm
L_X10Y70VDD_X10Y80VDD X10Y75VDD X10Y80VDD 2.91e-06nH
R_X10Y70VSS_X10Y80VSS X10Y70VSS X10Y75VSS 25mOhm
L_X10Y70VSS_X10Y80VSS X10Y75VSS X10Y80VSS 2.91e-06nH
R_X10Y80VDD_X10Y90VDD X10Y80VDD X10Y85VDD 25mOhm
L_X10Y80VDD_X10Y90VDD X10Y85VDD X10Y90VDD 2.91e-06nH
R_X10Y80VSS_X10Y90VSS X10Y80VSS X10Y85VSS 25mOhm
L_X10Y80VSS_X10Y90VSS X10Y85VSS X10Y90VSS 2.91e-06nH
R_X10Y90VDD_X10Y100VDD X10Y90VDD X10Y95VDD 25mOhm
L_X10Y90VDD_X10Y100VDD X10Y95VDD X10Y100VDD 2.91e-06nH
R_X10Y90VSS_X10Y100VSS X10Y90VSS X10Y95VSS 25mOhm
L_X10Y90VSS_X10Y100VSS X10Y95VSS X10Y100VSS 2.91e-06nH
R_X10Y100VDD_X10Y110VDD X10Y100VDD X10Y105VDD 25mOhm
L_X10Y100VDD_X10Y110VDD X10Y105VDD X10Y110VDD 2.91e-06nH
R_X10Y100VSS_X10Y110VSS X10Y100VSS X10Y105VSS 25mOhm
L_X10Y100VSS_X10Y110VSS X10Y105VSS X10Y110VSS 2.91e-06nH
R_X10Y110VDD_X10Y120VDD X10Y110VDD X10Y115VDD 25mOhm
L_X10Y110VDD_X10Y120VDD X10Y115VDD X10Y120VDD 2.91e-06nH
R_X10Y110VSS_X10Y120VSS X10Y110VSS X10Y115VSS 25mOhm
L_X10Y110VSS_X10Y120VSS X10Y115VSS X10Y120VSS 2.91e-06nH
R_X20Y10VDD_X20Y20VDD X20Y10VDD X20Y15VDD 25mOhm
L_X20Y10VDD_X20Y20VDD X20Y15VDD X20Y20VDD 2.91e-06nH
R_X20Y10VSS_X20Y20VSS X20Y10VSS X20Y15VSS 25mOhm
L_X20Y10VSS_X20Y20VSS X20Y15VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X20Y30VDD X20Y20VDD X20Y25VDD 25mOhm
L_X20Y20VDD_X20Y30VDD X20Y25VDD X20Y30VDD 2.91e-06nH
R_X20Y20VSS_X20Y30VSS X20Y20VSS X20Y25VSS 25mOhm
L_X20Y20VSS_X20Y30VSS X20Y25VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X20Y40VDD X20Y30VDD X20Y35VDD 25mOhm
L_X20Y30VDD_X20Y40VDD X20Y35VDD X20Y40VDD 2.91e-06nH
R_X20Y30VSS_X20Y40VSS X20Y30VSS X20Y35VSS 25mOhm
L_X20Y30VSS_X20Y40VSS X20Y35VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X20Y50VDD X20Y40VDD X20Y45VDD 25mOhm
L_X20Y40VDD_X20Y50VDD X20Y45VDD X20Y50VDD 2.91e-06nH
R_X20Y40VSS_X20Y50VSS X20Y40VSS X20Y45VSS 25mOhm
L_X20Y40VSS_X20Y50VSS X20Y45VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X20Y60VDD X20Y50VDD X20Y55VDD 25mOhm
L_X20Y50VDD_X20Y60VDD X20Y55VDD X20Y60VDD 2.91e-06nH
R_X20Y50VSS_X20Y60VSS X20Y50VSS X20Y55VSS 25mOhm
L_X20Y50VSS_X20Y60VSS X20Y55VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X20Y70VDD X20Y60VDD X20Y65VDD 25mOhm
L_X20Y60VDD_X20Y70VDD X20Y65VDD X20Y70VDD 2.91e-06nH
R_X20Y60VSS_X20Y70VSS X20Y60VSS X20Y65VSS 25mOhm
L_X20Y60VSS_X20Y70VSS X20Y65VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X20Y80VDD X20Y70VDD X20Y75VDD 25mOhm
L_X20Y70VDD_X20Y80VDD X20Y75VDD X20Y80VDD 2.91e-06nH
R_X20Y70VSS_X20Y80VSS X20Y70VSS X20Y75VSS 25mOhm
L_X20Y70VSS_X20Y80VSS X20Y75VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X20Y90VDD X20Y80VDD X20Y85VDD 25mOhm
L_X20Y80VDD_X20Y90VDD X20Y85VDD X20Y90VDD 2.91e-06nH
R_X20Y80VSS_X20Y90VSS X20Y80VSS X20Y85VSS 25mOhm
L_X20Y80VSS_X20Y90VSS X20Y85VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X20Y100VDD X20Y90VDD X20Y95VDD 25mOhm
L_X20Y90VDD_X20Y100VDD X20Y95VDD X20Y100VDD 2.91e-06nH
R_X20Y90VSS_X20Y100VSS X20Y90VSS X20Y95VSS 25mOhm
L_X20Y90VSS_X20Y100VSS X20Y95VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X20Y110VDD X20Y100VDD X20Y105VDD 25mOhm
L_X20Y100VDD_X20Y110VDD X20Y105VDD X20Y110VDD 2.91e-06nH
R_X20Y100VSS_X20Y110VSS X20Y100VSS X20Y105VSS 25mOhm
L_X20Y100VSS_X20Y110VSS X20Y105VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X20Y120VDD X20Y110VDD X20Y115VDD 25mOhm
L_X20Y110VDD_X20Y120VDD X20Y115VDD X20Y120VDD 2.91e-06nH
R_X20Y110VSS_X20Y120VSS X20Y110VSS X20Y115VSS 25mOhm
L_X20Y110VSS_X20Y120VSS X20Y115VSS X20Y120VSS 2.91e-06nH
R_X30Y10VDD_X30Y20VDD X30Y10VDD X30Y15VDD 25mOhm
L_X30Y10VDD_X30Y20VDD X30Y15VDD X30Y20VDD 2.91e-06nH
R_X30Y10VSS_X30Y20VSS X30Y10VSS X30Y15VSS 25mOhm
L_X30Y10VSS_X30Y20VSS X30Y15VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X30Y30VDD X30Y20VDD X30Y25VDD 25mOhm
L_X30Y20VDD_X30Y30VDD X30Y25VDD X30Y30VDD 2.91e-06nH
R_X30Y20VSS_X30Y30VSS X30Y20VSS X30Y25VSS 25mOhm
L_X30Y20VSS_X30Y30VSS X30Y25VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X30Y40VDD X30Y30VDD X30Y35VDD 25mOhm
L_X30Y30VDD_X30Y40VDD X30Y35VDD X30Y40VDD 2.91e-06nH
R_X30Y30VSS_X30Y40VSS X30Y30VSS X30Y35VSS 25mOhm
L_X30Y30VSS_X30Y40VSS X30Y35VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X30Y50VDD X30Y40VDD X30Y45VDD 25mOhm
L_X30Y40VDD_X30Y50VDD X30Y45VDD X30Y50VDD 2.91e-06nH
R_X30Y40VSS_X30Y50VSS X30Y40VSS X30Y45VSS 25mOhm
L_X30Y40VSS_X30Y50VSS X30Y45VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X30Y60VDD X30Y50VDD X30Y55VDD 25mOhm
L_X30Y50VDD_X30Y60VDD X30Y55VDD X30Y60VDD 2.91e-06nH
R_X30Y50VSS_X30Y60VSS X30Y50VSS X30Y55VSS 25mOhm
L_X30Y50VSS_X30Y60VSS X30Y55VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X30Y70VDD X30Y60VDD X30Y65VDD 25mOhm
L_X30Y60VDD_X30Y70VDD X30Y65VDD X30Y70VDD 2.91e-06nH
R_X30Y60VSS_X30Y70VSS X30Y60VSS X30Y65VSS 25mOhm
L_X30Y60VSS_X30Y70VSS X30Y65VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X30Y80VDD X30Y70VDD X30Y75VDD 25mOhm
L_X30Y70VDD_X30Y80VDD X30Y75VDD X30Y80VDD 2.91e-06nH
R_X30Y70VSS_X30Y80VSS X30Y70VSS X30Y75VSS 25mOhm
L_X30Y70VSS_X30Y80VSS X30Y75VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X30Y90VDD X30Y80VDD X30Y85VDD 25mOhm
L_X30Y80VDD_X30Y90VDD X30Y85VDD X30Y90VDD 2.91e-06nH
R_X30Y80VSS_X30Y90VSS X30Y80VSS X30Y85VSS 25mOhm
L_X30Y80VSS_X30Y90VSS X30Y85VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X30Y100VDD X30Y90VDD X30Y95VDD 25mOhm
L_X30Y90VDD_X30Y100VDD X30Y95VDD X30Y100VDD 2.91e-06nH
R_X30Y90VSS_X30Y100VSS X30Y90VSS X30Y95VSS 25mOhm
L_X30Y90VSS_X30Y100VSS X30Y95VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X30Y110VDD X30Y100VDD X30Y105VDD 25mOhm
L_X30Y100VDD_X30Y110VDD X30Y105VDD X30Y110VDD 2.91e-06nH
R_X30Y100VSS_X30Y110VSS X30Y100VSS X30Y105VSS 25mOhm
L_X30Y100VSS_X30Y110VSS X30Y105VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X30Y120VDD X30Y110VDD X30Y115VDD 25mOhm
L_X30Y110VDD_X30Y120VDD X30Y115VDD X30Y120VDD 2.91e-06nH
R_X30Y110VSS_X30Y120VSS X30Y110VSS X30Y115VSS 25mOhm
L_X30Y110VSS_X30Y120VSS X30Y115VSS X30Y120VSS 2.91e-06nH
R_X40Y10VDD_X40Y20VDD X40Y10VDD X40Y15VDD 25mOhm
L_X40Y10VDD_X40Y20VDD X40Y15VDD X40Y20VDD 2.91e-06nH
R_X40Y10VSS_X40Y20VSS X40Y10VSS X40Y15VSS 25mOhm
L_X40Y10VSS_X40Y20VSS X40Y15VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X40Y30VDD X40Y20VDD X40Y25VDD 25mOhm
L_X40Y20VDD_X40Y30VDD X40Y25VDD X40Y30VDD 2.91e-06nH
R_X40Y20VSS_X40Y30VSS X40Y20VSS X40Y25VSS 25mOhm
L_X40Y20VSS_X40Y30VSS X40Y25VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X40Y40VDD X40Y30VDD X40Y35VDD 25mOhm
L_X40Y30VDD_X40Y40VDD X40Y35VDD X40Y40VDD 2.91e-06nH
R_X40Y30VSS_X40Y40VSS X40Y30VSS X40Y35VSS 25mOhm
L_X40Y30VSS_X40Y40VSS X40Y35VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X40Y50VDD X40Y40VDD X40Y45VDD 25mOhm
L_X40Y40VDD_X40Y50VDD X40Y45VDD X40Y50VDD 2.91e-06nH
R_X40Y40VSS_X40Y50VSS X40Y40VSS X40Y45VSS 25mOhm
L_X40Y40VSS_X40Y50VSS X40Y45VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X40Y60VDD X40Y50VDD X40Y55VDD 25mOhm
L_X40Y50VDD_X40Y60VDD X40Y55VDD X40Y60VDD 2.91e-06nH
R_X40Y50VSS_X40Y60VSS X40Y50VSS X40Y55VSS 25mOhm
L_X40Y50VSS_X40Y60VSS X40Y55VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X40Y70VDD X40Y60VDD X40Y65VDD 25mOhm
L_X40Y60VDD_X40Y70VDD X40Y65VDD X40Y70VDD 2.91e-06nH
R_X40Y60VSS_X40Y70VSS X40Y60VSS X40Y65VSS 25mOhm
L_X40Y60VSS_X40Y70VSS X40Y65VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X40Y80VDD X40Y70VDD X40Y75VDD 25mOhm
L_X40Y70VDD_X40Y80VDD X40Y75VDD X40Y80VDD 2.91e-06nH
R_X40Y70VSS_X40Y80VSS X40Y70VSS X40Y75VSS 25mOhm
L_X40Y70VSS_X40Y80VSS X40Y75VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X40Y90VDD X40Y80VDD X40Y85VDD 25mOhm
L_X40Y80VDD_X40Y90VDD X40Y85VDD X40Y90VDD 2.91e-06nH
R_X40Y80VSS_X40Y90VSS X40Y80VSS X40Y85VSS 25mOhm
L_X40Y80VSS_X40Y90VSS X40Y85VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X40Y100VDD X40Y90VDD X40Y95VDD 25mOhm
L_X40Y90VDD_X40Y100VDD X40Y95VDD X40Y100VDD 2.91e-06nH
R_X40Y90VSS_X40Y100VSS X40Y90VSS X40Y95VSS 25mOhm
L_X40Y90VSS_X40Y100VSS X40Y95VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X40Y110VDD X40Y100VDD X40Y105VDD 25mOhm
L_X40Y100VDD_X40Y110VDD X40Y105VDD X40Y110VDD 2.91e-06nH
R_X40Y100VSS_X40Y110VSS X40Y100VSS X40Y105VSS 25mOhm
L_X40Y100VSS_X40Y110VSS X40Y105VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X40Y120VDD X40Y110VDD X40Y115VDD 25mOhm
L_X40Y110VDD_X40Y120VDD X40Y115VDD X40Y120VDD 2.91e-06nH
R_X40Y110VSS_X40Y120VSS X40Y110VSS X40Y115VSS 25mOhm
L_X40Y110VSS_X40Y120VSS X40Y115VSS X40Y120VSS 2.91e-06nH
R_X50Y10VDD_X50Y20VDD X50Y10VDD X50Y15VDD 25mOhm
L_X50Y10VDD_X50Y20VDD X50Y15VDD X50Y20VDD 2.91e-06nH
R_X50Y10VSS_X50Y20VSS X50Y10VSS X50Y15VSS 25mOhm
L_X50Y10VSS_X50Y20VSS X50Y15VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X50Y30VDD X50Y20VDD X50Y25VDD 25mOhm
L_X50Y20VDD_X50Y30VDD X50Y25VDD X50Y30VDD 2.91e-06nH
R_X50Y20VSS_X50Y30VSS X50Y20VSS X50Y25VSS 25mOhm
L_X50Y20VSS_X50Y30VSS X50Y25VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X50Y40VDD X50Y30VDD X50Y35VDD 25mOhm
L_X50Y30VDD_X50Y40VDD X50Y35VDD X50Y40VDD 2.91e-06nH
R_X50Y30VSS_X50Y40VSS X50Y30VSS X50Y35VSS 25mOhm
L_X50Y30VSS_X50Y40VSS X50Y35VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X50Y50VDD X50Y40VDD X50Y45VDD 25mOhm
L_X50Y40VDD_X50Y50VDD X50Y45VDD X50Y50VDD 2.91e-06nH
R_X50Y40VSS_X50Y50VSS X50Y40VSS X50Y45VSS 25mOhm
L_X50Y40VSS_X50Y50VSS X50Y45VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X50Y60VDD X50Y50VDD X50Y55VDD 25mOhm
L_X50Y50VDD_X50Y60VDD X50Y55VDD X50Y60VDD 2.91e-06nH
R_X50Y50VSS_X50Y60VSS X50Y50VSS X50Y55VSS 25mOhm
L_X50Y50VSS_X50Y60VSS X50Y55VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X50Y70VDD X50Y60VDD X50Y65VDD 25mOhm
L_X50Y60VDD_X50Y70VDD X50Y65VDD X50Y70VDD 2.91e-06nH
R_X50Y60VSS_X50Y70VSS X50Y60VSS X50Y65VSS 25mOhm
L_X50Y60VSS_X50Y70VSS X50Y65VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X50Y80VDD X50Y70VDD X50Y75VDD 25mOhm
L_X50Y70VDD_X50Y80VDD X50Y75VDD X50Y80VDD 2.91e-06nH
R_X50Y70VSS_X50Y80VSS X50Y70VSS X50Y75VSS 25mOhm
L_X50Y70VSS_X50Y80VSS X50Y75VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X50Y90VDD X50Y80VDD X50Y85VDD 25mOhm
L_X50Y80VDD_X50Y90VDD X50Y85VDD X50Y90VDD 2.91e-06nH
R_X50Y80VSS_X50Y90VSS X50Y80VSS X50Y85VSS 25mOhm
L_X50Y80VSS_X50Y90VSS X50Y85VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X50Y100VDD X50Y90VDD X50Y95VDD 25mOhm
L_X50Y90VDD_X50Y100VDD X50Y95VDD X50Y100VDD 2.91e-06nH
R_X50Y90VSS_X50Y100VSS X50Y90VSS X50Y95VSS 25mOhm
L_X50Y90VSS_X50Y100VSS X50Y95VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X50Y110VDD X50Y100VDD X50Y105VDD 25mOhm
L_X50Y100VDD_X50Y110VDD X50Y105VDD X50Y110VDD 2.91e-06nH
R_X50Y100VSS_X50Y110VSS X50Y100VSS X50Y105VSS 25mOhm
L_X50Y100VSS_X50Y110VSS X50Y105VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X50Y120VDD X50Y110VDD X50Y115VDD 25mOhm
L_X50Y110VDD_X50Y120VDD X50Y115VDD X50Y120VDD 2.91e-06nH
R_X50Y110VSS_X50Y120VSS X50Y110VSS X50Y115VSS 25mOhm
L_X50Y110VSS_X50Y120VSS X50Y115VSS X50Y120VSS 2.91e-06nH
R_X60Y10VDD_X60Y20VDD X60Y10VDD X60Y15VDD 25mOhm
L_X60Y10VDD_X60Y20VDD X60Y15VDD X60Y20VDD 2.91e-06nH
R_X60Y10VSS_X60Y20VSS X60Y10VSS X60Y15VSS 25mOhm
L_X60Y10VSS_X60Y20VSS X60Y15VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X60Y30VDD X60Y20VDD X60Y25VDD 25mOhm
L_X60Y20VDD_X60Y30VDD X60Y25VDD X60Y30VDD 2.91e-06nH
R_X60Y20VSS_X60Y30VSS X60Y20VSS X60Y25VSS 25mOhm
L_X60Y20VSS_X60Y30VSS X60Y25VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X60Y40VDD X60Y30VDD X60Y35VDD 25mOhm
L_X60Y30VDD_X60Y40VDD X60Y35VDD X60Y40VDD 2.91e-06nH
R_X60Y30VSS_X60Y40VSS X60Y30VSS X60Y35VSS 25mOhm
L_X60Y30VSS_X60Y40VSS X60Y35VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X60Y50VDD X60Y40VDD X60Y45VDD 25mOhm
L_X60Y40VDD_X60Y50VDD X60Y45VDD X60Y50VDD 2.91e-06nH
R_X60Y40VSS_X60Y50VSS X60Y40VSS X60Y45VSS 25mOhm
L_X60Y40VSS_X60Y50VSS X60Y45VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X60Y60VDD X60Y50VDD X60Y55VDD 25mOhm
L_X60Y50VDD_X60Y60VDD X60Y55VDD X60Y60VDD 2.91e-06nH
R_X60Y50VSS_X60Y60VSS X60Y50VSS X60Y55VSS 25mOhm
L_X60Y50VSS_X60Y60VSS X60Y55VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X60Y70VDD X60Y60VDD X60Y65VDD 25mOhm
L_X60Y60VDD_X60Y70VDD X60Y65VDD X60Y70VDD 2.91e-06nH
R_X60Y60VSS_X60Y70VSS X60Y60VSS X60Y65VSS 25mOhm
L_X60Y60VSS_X60Y70VSS X60Y65VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X60Y80VDD X60Y70VDD X60Y75VDD 25mOhm
L_X60Y70VDD_X60Y80VDD X60Y75VDD X60Y80VDD 2.91e-06nH
R_X60Y70VSS_X60Y80VSS X60Y70VSS X60Y75VSS 25mOhm
L_X60Y70VSS_X60Y80VSS X60Y75VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X60Y90VDD X60Y80VDD X60Y85VDD 25mOhm
L_X60Y80VDD_X60Y90VDD X60Y85VDD X60Y90VDD 2.91e-06nH
R_X60Y80VSS_X60Y90VSS X60Y80VSS X60Y85VSS 25mOhm
L_X60Y80VSS_X60Y90VSS X60Y85VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X60Y100VDD X60Y90VDD X60Y95VDD 25mOhm
L_X60Y90VDD_X60Y100VDD X60Y95VDD X60Y100VDD 2.91e-06nH
R_X60Y90VSS_X60Y100VSS X60Y90VSS X60Y95VSS 25mOhm
L_X60Y90VSS_X60Y100VSS X60Y95VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X60Y110VDD X60Y100VDD X60Y105VDD 25mOhm
L_X60Y100VDD_X60Y110VDD X60Y105VDD X60Y110VDD 2.91e-06nH
R_X60Y100VSS_X60Y110VSS X60Y100VSS X60Y105VSS 25mOhm
L_X60Y100VSS_X60Y110VSS X60Y105VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X60Y120VDD X60Y110VDD X60Y115VDD 25mOhm
L_X60Y110VDD_X60Y120VDD X60Y115VDD X60Y120VDD 2.91e-06nH
R_X60Y110VSS_X60Y120VSS X60Y110VSS X60Y115VSS 25mOhm
L_X60Y110VSS_X60Y120VSS X60Y115VSS X60Y120VSS 2.91e-06nH
R_X70Y10VDD_X70Y20VDD X70Y10VDD X70Y15VDD 25mOhm
L_X70Y10VDD_X70Y20VDD X70Y15VDD X70Y20VDD 2.91e-06nH
R_X70Y10VSS_X70Y20VSS X70Y10VSS X70Y15VSS 25mOhm
L_X70Y10VSS_X70Y20VSS X70Y15VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X70Y30VDD X70Y20VDD X70Y25VDD 25mOhm
L_X70Y20VDD_X70Y30VDD X70Y25VDD X70Y30VDD 2.91e-06nH
R_X70Y20VSS_X70Y30VSS X70Y20VSS X70Y25VSS 25mOhm
L_X70Y20VSS_X70Y30VSS X70Y25VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X70Y40VDD X70Y30VDD X70Y35VDD 25mOhm
L_X70Y30VDD_X70Y40VDD X70Y35VDD X70Y40VDD 2.91e-06nH
R_X70Y30VSS_X70Y40VSS X70Y30VSS X70Y35VSS 25mOhm
L_X70Y30VSS_X70Y40VSS X70Y35VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X70Y50VDD X70Y40VDD X70Y45VDD 25mOhm
L_X70Y40VDD_X70Y50VDD X70Y45VDD X70Y50VDD 2.91e-06nH
R_X70Y40VSS_X70Y50VSS X70Y40VSS X70Y45VSS 25mOhm
L_X70Y40VSS_X70Y50VSS X70Y45VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X70Y60VDD X70Y50VDD X70Y55VDD 25mOhm
L_X70Y50VDD_X70Y60VDD X70Y55VDD X70Y60VDD 2.91e-06nH
R_X70Y50VSS_X70Y60VSS X70Y50VSS X70Y55VSS 25mOhm
L_X70Y50VSS_X70Y60VSS X70Y55VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X70Y70VDD X70Y60VDD X70Y65VDD 25mOhm
L_X70Y60VDD_X70Y70VDD X70Y65VDD X70Y70VDD 2.91e-06nH
R_X70Y60VSS_X70Y70VSS X70Y60VSS X70Y65VSS 25mOhm
L_X70Y60VSS_X70Y70VSS X70Y65VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X70Y80VDD X70Y70VDD X70Y75VDD 25mOhm
L_X70Y70VDD_X70Y80VDD X70Y75VDD X70Y80VDD 2.91e-06nH
R_X70Y70VSS_X70Y80VSS X70Y70VSS X70Y75VSS 25mOhm
L_X70Y70VSS_X70Y80VSS X70Y75VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X70Y90VDD X70Y80VDD X70Y85VDD 25mOhm
L_X70Y80VDD_X70Y90VDD X70Y85VDD X70Y90VDD 2.91e-06nH
R_X70Y80VSS_X70Y90VSS X70Y80VSS X70Y85VSS 25mOhm
L_X70Y80VSS_X70Y90VSS X70Y85VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X70Y100VDD X70Y90VDD X70Y95VDD 25mOhm
L_X70Y90VDD_X70Y100VDD X70Y95VDD X70Y100VDD 2.91e-06nH
R_X70Y90VSS_X70Y100VSS X70Y90VSS X70Y95VSS 25mOhm
L_X70Y90VSS_X70Y100VSS X70Y95VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X70Y110VDD X70Y100VDD X70Y105VDD 25mOhm
L_X70Y100VDD_X70Y110VDD X70Y105VDD X70Y110VDD 2.91e-06nH
R_X70Y100VSS_X70Y110VSS X70Y100VSS X70Y105VSS 25mOhm
L_X70Y100VSS_X70Y110VSS X70Y105VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X70Y120VDD X70Y110VDD X70Y115VDD 25mOhm
L_X70Y110VDD_X70Y120VDD X70Y115VDD X70Y120VDD 2.91e-06nH
R_X70Y110VSS_X70Y120VSS X70Y110VSS X70Y115VSS 25mOhm
L_X70Y110VSS_X70Y120VSS X70Y115VSS X70Y120VSS 2.91e-06nH
R_X80Y10VDD_X80Y20VDD X80Y10VDD X80Y15VDD 25mOhm
L_X80Y10VDD_X80Y20VDD X80Y15VDD X80Y20VDD 2.91e-06nH
R_X80Y10VSS_X80Y20VSS X80Y10VSS X80Y15VSS 25mOhm
L_X80Y10VSS_X80Y20VSS X80Y15VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X80Y30VDD X80Y20VDD X80Y25VDD 25mOhm
L_X80Y20VDD_X80Y30VDD X80Y25VDD X80Y30VDD 2.91e-06nH
R_X80Y20VSS_X80Y30VSS X80Y20VSS X80Y25VSS 25mOhm
L_X80Y20VSS_X80Y30VSS X80Y25VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X80Y40VDD X80Y30VDD X80Y35VDD 25mOhm
L_X80Y30VDD_X80Y40VDD X80Y35VDD X80Y40VDD 2.91e-06nH
R_X80Y30VSS_X80Y40VSS X80Y30VSS X80Y35VSS 25mOhm
L_X80Y30VSS_X80Y40VSS X80Y35VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X80Y50VDD X80Y40VDD X80Y45VDD 25mOhm
L_X80Y40VDD_X80Y50VDD X80Y45VDD X80Y50VDD 2.91e-06nH
R_X80Y40VSS_X80Y50VSS X80Y40VSS X80Y45VSS 25mOhm
L_X80Y40VSS_X80Y50VSS X80Y45VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X80Y60VDD X80Y50VDD X80Y55VDD 25mOhm
L_X80Y50VDD_X80Y60VDD X80Y55VDD X80Y60VDD 2.91e-06nH
R_X80Y50VSS_X80Y60VSS X80Y50VSS X80Y55VSS 25mOhm
L_X80Y50VSS_X80Y60VSS X80Y55VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X80Y70VDD X80Y60VDD X80Y65VDD 25mOhm
L_X80Y60VDD_X80Y70VDD X80Y65VDD X80Y70VDD 2.91e-06nH
R_X80Y60VSS_X80Y70VSS X80Y60VSS X80Y65VSS 25mOhm
L_X80Y60VSS_X80Y70VSS X80Y65VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X80Y80VDD X80Y70VDD X80Y75VDD 25mOhm
L_X80Y70VDD_X80Y80VDD X80Y75VDD X80Y80VDD 2.91e-06nH
R_X80Y70VSS_X80Y80VSS X80Y70VSS X80Y75VSS 25mOhm
L_X80Y70VSS_X80Y80VSS X80Y75VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X80Y90VDD X80Y80VDD X80Y85VDD 25mOhm
L_X80Y80VDD_X80Y90VDD X80Y85VDD X80Y90VDD 2.91e-06nH
R_X80Y80VSS_X80Y90VSS X80Y80VSS X80Y85VSS 25mOhm
L_X80Y80VSS_X80Y90VSS X80Y85VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X80Y100VDD X80Y90VDD X80Y95VDD 25mOhm
L_X80Y90VDD_X80Y100VDD X80Y95VDD X80Y100VDD 2.91e-06nH
R_X80Y90VSS_X80Y100VSS X80Y90VSS X80Y95VSS 25mOhm
L_X80Y90VSS_X80Y100VSS X80Y95VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X80Y110VDD X80Y100VDD X80Y105VDD 25mOhm
L_X80Y100VDD_X80Y110VDD X80Y105VDD X80Y110VDD 2.91e-06nH
R_X80Y100VSS_X80Y110VSS X80Y100VSS X80Y105VSS 25mOhm
L_X80Y100VSS_X80Y110VSS X80Y105VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X80Y120VDD X80Y110VDD X80Y115VDD 25mOhm
L_X80Y110VDD_X80Y120VDD X80Y115VDD X80Y120VDD 2.91e-06nH
R_X80Y110VSS_X80Y120VSS X80Y110VSS X80Y115VSS 25mOhm
L_X80Y110VSS_X80Y120VSS X80Y115VSS X80Y120VSS 2.91e-06nH
R_X90Y10VDD_X90Y20VDD X90Y10VDD X90Y15VDD 25mOhm
L_X90Y10VDD_X90Y20VDD X90Y15VDD X90Y20VDD 2.91e-06nH
R_X90Y10VSS_X90Y20VSS X90Y10VSS X90Y15VSS 25mOhm
L_X90Y10VSS_X90Y20VSS X90Y15VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X90Y30VDD X90Y20VDD X90Y25VDD 25mOhm
L_X90Y20VDD_X90Y30VDD X90Y25VDD X90Y30VDD 2.91e-06nH
R_X90Y20VSS_X90Y30VSS X90Y20VSS X90Y25VSS 25mOhm
L_X90Y20VSS_X90Y30VSS X90Y25VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X90Y40VDD X90Y30VDD X90Y35VDD 25mOhm
L_X90Y30VDD_X90Y40VDD X90Y35VDD X90Y40VDD 2.91e-06nH
R_X90Y30VSS_X90Y40VSS X90Y30VSS X90Y35VSS 25mOhm
L_X90Y30VSS_X90Y40VSS X90Y35VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X90Y50VDD X90Y40VDD X90Y45VDD 25mOhm
L_X90Y40VDD_X90Y50VDD X90Y45VDD X90Y50VDD 2.91e-06nH
R_X90Y40VSS_X90Y50VSS X90Y40VSS X90Y45VSS 25mOhm
L_X90Y40VSS_X90Y50VSS X90Y45VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X90Y60VDD X90Y50VDD X90Y55VDD 25mOhm
L_X90Y50VDD_X90Y60VDD X90Y55VDD X90Y60VDD 2.91e-06nH
R_X90Y50VSS_X90Y60VSS X90Y50VSS X90Y55VSS 25mOhm
L_X90Y50VSS_X90Y60VSS X90Y55VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X90Y70VDD X90Y60VDD X90Y65VDD 25mOhm
L_X90Y60VDD_X90Y70VDD X90Y65VDD X90Y70VDD 2.91e-06nH
R_X90Y60VSS_X90Y70VSS X90Y60VSS X90Y65VSS 25mOhm
L_X90Y60VSS_X90Y70VSS X90Y65VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X90Y80VDD X90Y70VDD X90Y75VDD 25mOhm
L_X90Y70VDD_X90Y80VDD X90Y75VDD X90Y80VDD 2.91e-06nH
R_X90Y70VSS_X90Y80VSS X90Y70VSS X90Y75VSS 25mOhm
L_X90Y70VSS_X90Y80VSS X90Y75VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X90Y90VDD X90Y80VDD X90Y85VDD 25mOhm
L_X90Y80VDD_X90Y90VDD X90Y85VDD X90Y90VDD 2.91e-06nH
R_X90Y80VSS_X90Y90VSS X90Y80VSS X90Y85VSS 25mOhm
L_X90Y80VSS_X90Y90VSS X90Y85VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X90Y100VDD X90Y90VDD X90Y95VDD 25mOhm
L_X90Y90VDD_X90Y100VDD X90Y95VDD X90Y100VDD 2.91e-06nH
R_X90Y90VSS_X90Y100VSS X90Y90VSS X90Y95VSS 25mOhm
L_X90Y90VSS_X90Y100VSS X90Y95VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X90Y110VDD X90Y100VDD X90Y105VDD 25mOhm
L_X90Y100VDD_X90Y110VDD X90Y105VDD X90Y110VDD 2.91e-06nH
R_X90Y100VSS_X90Y110VSS X90Y100VSS X90Y105VSS 25mOhm
L_X90Y100VSS_X90Y110VSS X90Y105VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X90Y120VDD X90Y110VDD X90Y115VDD 25mOhm
L_X90Y110VDD_X90Y120VDD X90Y115VDD X90Y120VDD 2.91e-06nH
R_X90Y110VSS_X90Y120VSS X90Y110VSS X90Y115VSS 25mOhm
L_X90Y110VSS_X90Y120VSS X90Y115VSS X90Y120VSS 2.91e-06nH
R_X100Y10VDD_X100Y20VDD X100Y10VDD X100Y15VDD 25mOhm
L_X100Y10VDD_X100Y20VDD X100Y15VDD X100Y20VDD 2.91e-06nH
R_X100Y10VSS_X100Y20VSS X100Y10VSS X100Y15VSS 25mOhm
L_X100Y10VSS_X100Y20VSS X100Y15VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X100Y30VDD X100Y20VDD X100Y25VDD 25mOhm
L_X100Y20VDD_X100Y30VDD X100Y25VDD X100Y30VDD 2.91e-06nH
R_X100Y20VSS_X100Y30VSS X100Y20VSS X100Y25VSS 25mOhm
L_X100Y20VSS_X100Y30VSS X100Y25VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X100Y40VDD X100Y30VDD X100Y35VDD 25mOhm
L_X100Y30VDD_X100Y40VDD X100Y35VDD X100Y40VDD 2.91e-06nH
R_X100Y30VSS_X100Y40VSS X100Y30VSS X100Y35VSS 25mOhm
L_X100Y30VSS_X100Y40VSS X100Y35VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X100Y50VDD X100Y40VDD X100Y45VDD 25mOhm
L_X100Y40VDD_X100Y50VDD X100Y45VDD X100Y50VDD 2.91e-06nH
R_X100Y40VSS_X100Y50VSS X100Y40VSS X100Y45VSS 25mOhm
L_X100Y40VSS_X100Y50VSS X100Y45VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X100Y60VDD X100Y50VDD X100Y55VDD 25mOhm
L_X100Y50VDD_X100Y60VDD X100Y55VDD X100Y60VDD 2.91e-06nH
R_X100Y50VSS_X100Y60VSS X100Y50VSS X100Y55VSS 25mOhm
L_X100Y50VSS_X100Y60VSS X100Y55VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X100Y70VDD X100Y60VDD X100Y65VDD 25mOhm
L_X100Y60VDD_X100Y70VDD X100Y65VDD X100Y70VDD 2.91e-06nH
R_X100Y60VSS_X100Y70VSS X100Y60VSS X100Y65VSS 25mOhm
L_X100Y60VSS_X100Y70VSS X100Y65VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X100Y80VDD X100Y70VDD X100Y75VDD 25mOhm
L_X100Y70VDD_X100Y80VDD X100Y75VDD X100Y80VDD 2.91e-06nH
R_X100Y70VSS_X100Y80VSS X100Y70VSS X100Y75VSS 25mOhm
L_X100Y70VSS_X100Y80VSS X100Y75VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X100Y90VDD X100Y80VDD X100Y85VDD 25mOhm
L_X100Y80VDD_X100Y90VDD X100Y85VDD X100Y90VDD 2.91e-06nH
R_X100Y80VSS_X100Y90VSS X100Y80VSS X100Y85VSS 25mOhm
L_X100Y80VSS_X100Y90VSS X100Y85VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X100Y100VDD X100Y90VDD X100Y95VDD 25mOhm
L_X100Y90VDD_X100Y100VDD X100Y95VDD X100Y100VDD 2.91e-06nH
R_X100Y90VSS_X100Y100VSS X100Y90VSS X100Y95VSS 25mOhm
L_X100Y90VSS_X100Y100VSS X100Y95VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X100Y110VDD X100Y100VDD X100Y105VDD 25mOhm
L_X100Y100VDD_X100Y110VDD X100Y105VDD X100Y110VDD 2.91e-06nH
R_X100Y100VSS_X100Y110VSS X100Y100VSS X100Y105VSS 25mOhm
L_X100Y100VSS_X100Y110VSS X100Y105VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X100Y120VDD X100Y110VDD X100Y115VDD 25mOhm
L_X100Y110VDD_X100Y120VDD X100Y115VDD X100Y120VDD 2.91e-06nH
R_X100Y110VSS_X100Y120VSS X100Y110VSS X100Y115VSS 25mOhm
L_X100Y110VSS_X100Y120VSS X100Y115VSS X100Y120VSS 2.91e-06nH
R_X110Y10VDD_X110Y20VDD X110Y10VDD X110Y15VDD 25mOhm
L_X110Y10VDD_X110Y20VDD X110Y15VDD X110Y20VDD 2.91e-06nH
R_X110Y10VSS_X110Y20VSS X110Y10VSS X110Y15VSS 25mOhm
L_X110Y10VSS_X110Y20VSS X110Y15VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X110Y30VDD X110Y20VDD X110Y25VDD 25mOhm
L_X110Y20VDD_X110Y30VDD X110Y25VDD X110Y30VDD 2.91e-06nH
R_X110Y20VSS_X110Y30VSS X110Y20VSS X110Y25VSS 25mOhm
L_X110Y20VSS_X110Y30VSS X110Y25VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X110Y40VDD X110Y30VDD X110Y35VDD 25mOhm
L_X110Y30VDD_X110Y40VDD X110Y35VDD X110Y40VDD 2.91e-06nH
R_X110Y30VSS_X110Y40VSS X110Y30VSS X110Y35VSS 25mOhm
L_X110Y30VSS_X110Y40VSS X110Y35VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X110Y50VDD X110Y40VDD X110Y45VDD 25mOhm
L_X110Y40VDD_X110Y50VDD X110Y45VDD X110Y50VDD 2.91e-06nH
R_X110Y40VSS_X110Y50VSS X110Y40VSS X110Y45VSS 25mOhm
L_X110Y40VSS_X110Y50VSS X110Y45VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X110Y60VDD X110Y50VDD X110Y55VDD 25mOhm
L_X110Y50VDD_X110Y60VDD X110Y55VDD X110Y60VDD 2.91e-06nH
R_X110Y50VSS_X110Y60VSS X110Y50VSS X110Y55VSS 25mOhm
L_X110Y50VSS_X110Y60VSS X110Y55VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X110Y70VDD X110Y60VDD X110Y65VDD 25mOhm
L_X110Y60VDD_X110Y70VDD X110Y65VDD X110Y70VDD 2.91e-06nH
R_X110Y60VSS_X110Y70VSS X110Y60VSS X110Y65VSS 25mOhm
L_X110Y60VSS_X110Y70VSS X110Y65VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X110Y80VDD X110Y70VDD X110Y75VDD 25mOhm
L_X110Y70VDD_X110Y80VDD X110Y75VDD X110Y80VDD 2.91e-06nH
R_X110Y70VSS_X110Y80VSS X110Y70VSS X110Y75VSS 25mOhm
L_X110Y70VSS_X110Y80VSS X110Y75VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X110Y90VDD X110Y80VDD X110Y85VDD 25mOhm
L_X110Y80VDD_X110Y90VDD X110Y85VDD X110Y90VDD 2.91e-06nH
R_X110Y80VSS_X110Y90VSS X110Y80VSS X110Y85VSS 25mOhm
L_X110Y80VSS_X110Y90VSS X110Y85VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X110Y100VDD X110Y90VDD X110Y95VDD 25mOhm
L_X110Y90VDD_X110Y100VDD X110Y95VDD X110Y100VDD 2.91e-06nH
R_X110Y90VSS_X110Y100VSS X110Y90VSS X110Y95VSS 25mOhm
L_X110Y90VSS_X110Y100VSS X110Y95VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X110Y110VDD X110Y100VDD X110Y105VDD 25mOhm
L_X110Y100VDD_X110Y110VDD X110Y105VDD X110Y110VDD 2.91e-06nH
R_X110Y100VSS_X110Y110VSS X110Y100VSS X110Y105VSS 25mOhm
L_X110Y100VSS_X110Y110VSS X110Y105VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X110Y120VDD X110Y110VDD X110Y115VDD 25mOhm
L_X110Y110VDD_X110Y120VDD X110Y115VDD X110Y120VDD 2.91e-06nH
R_X110Y110VSS_X110Y120VSS X110Y110VSS X110Y115VSS 25mOhm
L_X110Y110VSS_X110Y120VSS X110Y115VSS X110Y120VSS 2.91e-06nH
R_X120Y10VDD_X120Y20VDD X120Y10VDD X120Y15VDD 25mOhm
L_X120Y10VDD_X120Y20VDD X120Y15VDD X120Y20VDD 2.91e-06nH
R_X120Y10VSS_X120Y20VSS X120Y10VSS X120Y15VSS 25mOhm
L_X120Y10VSS_X120Y20VSS X120Y15VSS X120Y20VSS 2.91e-06nH
R_X120Y20VDD_X120Y30VDD X120Y20VDD X120Y25VDD 25mOhm
L_X120Y20VDD_X120Y30VDD X120Y25VDD X120Y30VDD 2.91e-06nH
R_X120Y20VSS_X120Y30VSS X120Y20VSS X120Y25VSS 25mOhm
L_X120Y20VSS_X120Y30VSS X120Y25VSS X120Y30VSS 2.91e-06nH
R_X120Y30VDD_X120Y40VDD X120Y30VDD X120Y35VDD 25mOhm
L_X120Y30VDD_X120Y40VDD X120Y35VDD X120Y40VDD 2.91e-06nH
R_X120Y30VSS_X120Y40VSS X120Y30VSS X120Y35VSS 25mOhm
L_X120Y30VSS_X120Y40VSS X120Y35VSS X120Y40VSS 2.91e-06nH
R_X120Y40VDD_X120Y50VDD X120Y40VDD X120Y45VDD 25mOhm
L_X120Y40VDD_X120Y50VDD X120Y45VDD X120Y50VDD 2.91e-06nH
R_X120Y40VSS_X120Y50VSS X120Y40VSS X120Y45VSS 25mOhm
L_X120Y40VSS_X120Y50VSS X120Y45VSS X120Y50VSS 2.91e-06nH
R_X120Y50VDD_X120Y60VDD X120Y50VDD X120Y55VDD 25mOhm
L_X120Y50VDD_X120Y60VDD X120Y55VDD X120Y60VDD 2.91e-06nH
R_X120Y50VSS_X120Y60VSS X120Y50VSS X120Y55VSS 25mOhm
L_X120Y50VSS_X120Y60VSS X120Y55VSS X120Y60VSS 2.91e-06nH
R_X120Y60VDD_X120Y70VDD X120Y60VDD X120Y65VDD 25mOhm
L_X120Y60VDD_X120Y70VDD X120Y65VDD X120Y70VDD 2.91e-06nH
R_X120Y60VSS_X120Y70VSS X120Y60VSS X120Y65VSS 25mOhm
L_X120Y60VSS_X120Y70VSS X120Y65VSS X120Y70VSS 2.91e-06nH
R_X120Y70VDD_X120Y80VDD X120Y70VDD X120Y75VDD 25mOhm
L_X120Y70VDD_X120Y80VDD X120Y75VDD X120Y80VDD 2.91e-06nH
R_X120Y70VSS_X120Y80VSS X120Y70VSS X120Y75VSS 25mOhm
L_X120Y70VSS_X120Y80VSS X120Y75VSS X120Y80VSS 2.91e-06nH
R_X120Y80VDD_X120Y90VDD X120Y80VDD X120Y85VDD 25mOhm
L_X120Y80VDD_X120Y90VDD X120Y85VDD X120Y90VDD 2.91e-06nH
R_X120Y80VSS_X120Y90VSS X120Y80VSS X120Y85VSS 25mOhm
L_X120Y80VSS_X120Y90VSS X120Y85VSS X120Y90VSS 2.91e-06nH
R_X120Y90VDD_X120Y100VDD X120Y90VDD X120Y95VDD 25mOhm
L_X120Y90VDD_X120Y100VDD X120Y95VDD X120Y100VDD 2.91e-06nH
R_X120Y90VSS_X120Y100VSS X120Y90VSS X120Y95VSS 25mOhm
L_X120Y90VSS_X120Y100VSS X120Y95VSS X120Y100VSS 2.91e-06nH
R_X120Y100VDD_X120Y110VDD X120Y100VDD X120Y105VDD 25mOhm
L_X120Y100VDD_X120Y110VDD X120Y105VDD X120Y110VDD 2.91e-06nH
R_X120Y100VSS_X120Y110VSS X120Y100VSS X120Y105VSS 25mOhm
L_X120Y100VSS_X120Y110VSS X120Y105VSS X120Y110VSS 2.91e-06nH
R_X120Y110VDD_X120Y120VDD X120Y110VDD X120Y115VDD 25mOhm
L_X120Y110VDD_X120Y120VDD X120Y115VDD X120Y120VDD 2.91e-06nH
R_X120Y110VSS_X120Y120VSS X120Y110VSS X120Y115VSS 25mOhm
L_X120Y110VSS_X120Y120VSS X120Y115VSS X120Y120VSS 2.91e-06nH
C_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VSS 10nF
C_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VSS 10nF
C_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VSS 10nF
C_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VSS 10nF
C_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VSS 10nF
C_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VSS 10nF
C_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VSS 10nF
C_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VSS 10nF
C_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VSS 10nF
C_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VSS 10nF
C_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VSS 10nF
C_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VSS 10nF
C_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VSS 10nF
C_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VSS 10nF
C_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VSS 10nF
C_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VSS 10nF
C_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VSS 10nF
C_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VSS 10nF
C_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VSS 10nF
C_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VSS 10nF
C_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VSS 10nF
C_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VSS 10nF
C_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VSS 10nF
C_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VSS 10nF
C_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VSS 10nF
C_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VSS 10nF
C_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VSS 10nF
C_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VSS 10nF
C_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VSS 10nF
C_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VSS 10nF
C_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VSS 10nF
C_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VSS 10nF
C_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VSS 10nF
C_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VSS 10nF
C_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VSS 10nF
C_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VSS 10nF
C_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VSS 10nF
C_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VSS 10nF
C_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VSS 10nF
C_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VSS 10nF
C_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VSS 10nF
C_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VSS 10nF
C_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VSS 10nF
C_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VSS 10nF
C_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VSS 10nF
C_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VSS 10nF
C_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VSS 10nF
C_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VSS 10nF
C_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VSS 10nF
C_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VSS 10nF
C_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VSS 10nF
C_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VSS 10nF
C_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VSS 10nF
C_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VSS 10nF
C_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VSS 10nF
C_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VSS 10nF
C_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VSS 10nF
C_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VSS 10nF
C_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VSS 10nF
C_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VSS 10nF
C_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VSS 10nF
C_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VSS 10nF
C_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VSS 10nF
C_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VSS 10nF
C_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VSS 10nF
C_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VSS 10nF
C_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VSS 10nF
C_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VSS 10nF
C_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VSS 10nF
C_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VSS 10nF
C_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VSS 10nF
C_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VSS 10nF
C_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VSS 10nF
C_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VSS 10nF
C_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VSS 10nF
C_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VSS 10nF
C_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VSS 10nF
C_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VSS 10nF
C_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VSS 10nF
C_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VSS 10nF
C_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VSS 10nF
C_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VSS 10nF
C_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VSS 10nF
C_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VSS 10nF
C_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VSS 10nF
C_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VSS 10nF
C_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VSS 10nF
C_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VSS 10nF
C_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VSS 10nF
C_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VSS 10nF
C_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VSS 10nF
C_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VSS 10nF
C_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VSS 10nF
C_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VSS 10nF
C_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VSS 10nF
C_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VSS 10nF
C_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VSS 10nF
C_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VSS 10nF
C_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VSS 10nF
C_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VSS 10nF
C_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VSS 10nF
C_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VSS 10nF
C_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VSS 10nF
C_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VSS 10nF
C_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VSS 10nF
C_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VSS 10nF
C_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VSS 10nF
C_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VSS 10nF
C_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VSS 10nF
C_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VSS 10nF
C_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VSS 10nF
C_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VSS 10nF
C_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VSS 10nF
C_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VSS 10nF
C_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VSS 10nF
C_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VSS 10nF
C_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VSS 10nF
C_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VSS 10nF
C_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VSS 10nF
C_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VSS 10nF
C_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VSS 10nF
C_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VSS 10nF
C_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VSS 10nF
C_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VSS 10nF
C_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VSS 10nF
C_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VSS 10nF
C_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VSS 10nF
C_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VSS 10nF
C_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VSS 10nF
C_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VSS 10nF
C_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VSS 10nF
C_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VSS 10nF
C_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VSS 10nF
C_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VSS 10nF
C_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VSS 10nF
C_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VSS 10nF
C_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VSS 10nF
C_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VSS 10nF
C_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VSS 10nF
C_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VSS 10nF
C_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VSS 10nF
C_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VSS 10nF
C_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VSS 10nF
C_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VSS 10nF
I_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VDDDM 1 AC=0.006944444444444444
V_X120Y120VDD_X120Y120VSS X120Y120VDDDM X120Y120VSS 0
I_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VDDDM 1 AC=0.006944444444444444
V_X120Y10VDD_X120Y10VSS X120Y10VDDDM X120Y10VSS 0
I_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VDDDM 1 AC=0.006944444444444444
V_X120Y20VDD_X120Y20VSS X120Y20VDDDM X120Y20VSS 0
I_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VDDDM 1 AC=0.006944444444444444
V_X120Y30VDD_X120Y30VSS X120Y30VDDDM X120Y30VSS 0
I_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VDDDM 1 AC=0.006944444444444444
V_X120Y40VDD_X120Y40VSS X120Y40VDDDM X120Y40VSS 0
I_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VDDDM 1 AC=0.006944444444444444
V_X120Y50VDD_X120Y50VSS X120Y50VDDDM X120Y50VSS 0
I_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VDDDM 1 AC=0.006944444444444444
V_X120Y60VDD_X120Y60VSS X120Y60VDDDM X120Y60VSS 0
I_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VDDDM 1 AC=0.006944444444444444
V_X120Y70VDD_X120Y70VSS X120Y70VDDDM X120Y70VSS 0
I_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VDDDM 1 AC=0.006944444444444444
V_X120Y80VDD_X120Y80VSS X120Y80VDDDM X120Y80VSS 0
I_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VDDDM 1 AC=0.006944444444444444
V_X120Y90VDD_X120Y90VSS X120Y90VDDDM X120Y90VSS 0
I_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VDDDM 1 AC=0.006944444444444444
V_X120Y100VDD_X120Y100VSS X120Y100VDDDM X120Y100VSS 0
I_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VDDDM 1 AC=0.006944444444444444
V_X120Y110VDD_X120Y110VSS X120Y110VDDDM X120Y110VSS 0
I_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VDDDM 1 AC=0.006944444444444444
V_X10Y120VDD_X10Y120VSS X10Y120VDDDM X10Y120VSS 0
I_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VDDDM 1 AC=0.006944444444444444
V_X10Y10VDD_X10Y10VSS X10Y10VDDDM X10Y10VSS 0
I_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VDDDM 1 AC=0.006944444444444444
V_X10Y20VDD_X10Y20VSS X10Y20VDDDM X10Y20VSS 0
I_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VDDDM 1 AC=0.006944444444444444
V_X10Y30VDD_X10Y30VSS X10Y30VDDDM X10Y30VSS 0
I_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VDDDM 1 AC=0.006944444444444444
V_X10Y40VDD_X10Y40VSS X10Y40VDDDM X10Y40VSS 0
I_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VDDDM 1 AC=0.006944444444444444
V_X10Y50VDD_X10Y50VSS X10Y50VDDDM X10Y50VSS 0
I_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VDDDM 1 AC=0.006944444444444444
V_X10Y60VDD_X10Y60VSS X10Y60VDDDM X10Y60VSS 0
I_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VDDDM 1 AC=0.006944444444444444
V_X10Y70VDD_X10Y70VSS X10Y70VDDDM X10Y70VSS 0
I_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VDDDM 1 AC=0.006944444444444444
V_X10Y80VDD_X10Y80VSS X10Y80VDDDM X10Y80VSS 0
I_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VDDDM 1 AC=0.006944444444444444
V_X10Y90VDD_X10Y90VSS X10Y90VDDDM X10Y90VSS 0
I_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VDDDM 1 AC=0.006944444444444444
V_X10Y100VDD_X10Y100VSS X10Y100VDDDM X10Y100VSS 0
I_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VDDDM 1 AC=0.006944444444444444
V_X10Y110VDD_X10Y110VSS X10Y110VDDDM X10Y110VSS 0
I_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VDDDM 1 AC=0.006944444444444444
V_X20Y120VDD_X20Y120VSS X20Y120VDDDM X20Y120VSS 0
I_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VDDDM 1 AC=0.006944444444444444
V_X20Y10VDD_X20Y10VSS X20Y10VDDDM X20Y10VSS 0
I_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VDDDM 1 AC=0.006944444444444444
V_X20Y20VDD_X20Y20VSS X20Y20VDDDM X20Y20VSS 0
I_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VDDDM 1 AC=0.006944444444444444
V_X20Y30VDD_X20Y30VSS X20Y30VDDDM X20Y30VSS 0
I_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VDDDM 1 AC=0.006944444444444444
V_X20Y40VDD_X20Y40VSS X20Y40VDDDM X20Y40VSS 0
I_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VDDDM 1 AC=0.006944444444444444
V_X20Y50VDD_X20Y50VSS X20Y50VDDDM X20Y50VSS 0
I_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VDDDM 1 AC=0.006944444444444444
V_X20Y60VDD_X20Y60VSS X20Y60VDDDM X20Y60VSS 0
I_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VDDDM 1 AC=0.006944444444444444
V_X20Y70VDD_X20Y70VSS X20Y70VDDDM X20Y70VSS 0
I_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VDDDM 1 AC=0.006944444444444444
V_X20Y80VDD_X20Y80VSS X20Y80VDDDM X20Y80VSS 0
I_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VDDDM 1 AC=0.006944444444444444
V_X20Y90VDD_X20Y90VSS X20Y90VDDDM X20Y90VSS 0
I_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VDDDM 1 AC=0.006944444444444444
V_X20Y100VDD_X20Y100VSS X20Y100VDDDM X20Y100VSS 0
I_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VDDDM 1 AC=0.006944444444444444
V_X20Y110VDD_X20Y110VSS X20Y110VDDDM X20Y110VSS 0
I_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VDDDM 1 AC=0.006944444444444444
V_X30Y120VDD_X30Y120VSS X30Y120VDDDM X30Y120VSS 0
I_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VDDDM 1 AC=0.006944444444444444
V_X30Y10VDD_X30Y10VSS X30Y10VDDDM X30Y10VSS 0
I_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VDDDM 1 AC=0.006944444444444444
V_X30Y20VDD_X30Y20VSS X30Y20VDDDM X30Y20VSS 0
I_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VDDDM 1 AC=0.006944444444444444
V_X30Y30VDD_X30Y30VSS X30Y30VDDDM X30Y30VSS 0
I_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VDDDM 1 AC=0.006944444444444444
V_X30Y40VDD_X30Y40VSS X30Y40VDDDM X30Y40VSS 0
I_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VDDDM 1 AC=0.006944444444444444
V_X30Y50VDD_X30Y50VSS X30Y50VDDDM X30Y50VSS 0
I_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VDDDM 1 AC=0.006944444444444444
V_X30Y60VDD_X30Y60VSS X30Y60VDDDM X30Y60VSS 0
I_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VDDDM 1 AC=0.006944444444444444
V_X30Y70VDD_X30Y70VSS X30Y70VDDDM X30Y70VSS 0
I_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VDDDM 1 AC=0.006944444444444444
V_X30Y80VDD_X30Y80VSS X30Y80VDDDM X30Y80VSS 0
I_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VDDDM 1 AC=0.006944444444444444
V_X30Y90VDD_X30Y90VSS X30Y90VDDDM X30Y90VSS 0
I_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VDDDM 1 AC=0.006944444444444444
V_X30Y100VDD_X30Y100VSS X30Y100VDDDM X30Y100VSS 0
I_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VDDDM 1 AC=0.006944444444444444
V_X30Y110VDD_X30Y110VSS X30Y110VDDDM X30Y110VSS 0
I_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VDDDM 1 AC=0.006944444444444444
V_X40Y120VDD_X40Y120VSS X40Y120VDDDM X40Y120VSS 0
I_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VDDDM 1 AC=0.006944444444444444
V_X40Y10VDD_X40Y10VSS X40Y10VDDDM X40Y10VSS 0
I_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VDDDM 1 AC=0.006944444444444444
V_X40Y20VDD_X40Y20VSS X40Y20VDDDM X40Y20VSS 0
I_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VDDDM 1 AC=0.006944444444444444
V_X40Y30VDD_X40Y30VSS X40Y30VDDDM X40Y30VSS 0
I_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VDDDM 1 AC=0.006944444444444444
V_X40Y40VDD_X40Y40VSS X40Y40VDDDM X40Y40VSS 0
I_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VDDDM 1 AC=0.006944444444444444
V_X40Y50VDD_X40Y50VSS X40Y50VDDDM X40Y50VSS 0
I_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VDDDM 1 AC=0.006944444444444444
V_X40Y60VDD_X40Y60VSS X40Y60VDDDM X40Y60VSS 0
I_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VDDDM 1 AC=0.006944444444444444
V_X40Y70VDD_X40Y70VSS X40Y70VDDDM X40Y70VSS 0
I_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VDDDM 1 AC=0.006944444444444444
V_X40Y80VDD_X40Y80VSS X40Y80VDDDM X40Y80VSS 0
I_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VDDDM 1 AC=0.006944444444444444
V_X40Y90VDD_X40Y90VSS X40Y90VDDDM X40Y90VSS 0
I_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VDDDM 1 AC=0.006944444444444444
V_X40Y100VDD_X40Y100VSS X40Y100VDDDM X40Y100VSS 0
I_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VDDDM 1 AC=0.006944444444444444
V_X40Y110VDD_X40Y110VSS X40Y110VDDDM X40Y110VSS 0
I_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VDDDM 1 AC=0.006944444444444444
V_X50Y120VDD_X50Y120VSS X50Y120VDDDM X50Y120VSS 0
I_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VDDDM 1 AC=0.006944444444444444
V_X50Y10VDD_X50Y10VSS X50Y10VDDDM X50Y10VSS 0
I_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VDDDM 1 AC=0.006944444444444444
V_X50Y20VDD_X50Y20VSS X50Y20VDDDM X50Y20VSS 0
I_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VDDDM 1 AC=0.006944444444444444
V_X50Y30VDD_X50Y30VSS X50Y30VDDDM X50Y30VSS 0
I_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VDDDM 1 AC=0.006944444444444444
V_X50Y40VDD_X50Y40VSS X50Y40VDDDM X50Y40VSS 0
I_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VDDDM 1 AC=0.006944444444444444
V_X50Y50VDD_X50Y50VSS X50Y50VDDDM X50Y50VSS 0
I_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VDDDM 1 AC=0.006944444444444444
V_X50Y60VDD_X50Y60VSS X50Y60VDDDM X50Y60VSS 0
I_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VDDDM 1 AC=0.006944444444444444
V_X50Y70VDD_X50Y70VSS X50Y70VDDDM X50Y70VSS 0
I_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VDDDM 1 AC=0.006944444444444444
V_X50Y80VDD_X50Y80VSS X50Y80VDDDM X50Y80VSS 0
I_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VDDDM 1 AC=0.006944444444444444
V_X50Y90VDD_X50Y90VSS X50Y90VDDDM X50Y90VSS 0
I_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VDDDM 1 AC=0.006944444444444444
V_X50Y100VDD_X50Y100VSS X50Y100VDDDM X50Y100VSS 0
I_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VDDDM 1 AC=0.006944444444444444
V_X50Y110VDD_X50Y110VSS X50Y110VDDDM X50Y110VSS 0
I_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VDDDM 1 AC=0.006944444444444444
V_X60Y120VDD_X60Y120VSS X60Y120VDDDM X60Y120VSS 0
I_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VDDDM 1 AC=0.006944444444444444
V_X60Y10VDD_X60Y10VSS X60Y10VDDDM X60Y10VSS 0
I_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VDDDM 1 AC=0.006944444444444444
V_X60Y20VDD_X60Y20VSS X60Y20VDDDM X60Y20VSS 0
I_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VDDDM 1 AC=0.006944444444444444
V_X60Y30VDD_X60Y30VSS X60Y30VDDDM X60Y30VSS 0
I_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VDDDM 1 AC=0.006944444444444444
V_X60Y40VDD_X60Y40VSS X60Y40VDDDM X60Y40VSS 0
I_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VDDDM 1 AC=0.006944444444444444
V_X60Y50VDD_X60Y50VSS X60Y50VDDDM X60Y50VSS 0
I_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VDDDM 1 AC=0.006944444444444444
V_X60Y60VDD_X60Y60VSS X60Y60VDDDM X60Y60VSS 0
I_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VDDDM 1 AC=0.006944444444444444
V_X60Y70VDD_X60Y70VSS X60Y70VDDDM X60Y70VSS 0
I_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VDDDM 1 AC=0.006944444444444444
V_X60Y80VDD_X60Y80VSS X60Y80VDDDM X60Y80VSS 0
I_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VDDDM 1 AC=0.006944444444444444
V_X60Y90VDD_X60Y90VSS X60Y90VDDDM X60Y90VSS 0
I_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VDDDM 1 AC=0.006944444444444444
V_X60Y100VDD_X60Y100VSS X60Y100VDDDM X60Y100VSS 0
I_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VDDDM 1 AC=0.006944444444444444
V_X60Y110VDD_X60Y110VSS X60Y110VDDDM X60Y110VSS 0
I_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VDDDM 1 AC=0.006944444444444444
V_X70Y120VDD_X70Y120VSS X70Y120VDDDM X70Y120VSS 0
I_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VDDDM 1 AC=0.006944444444444444
V_X70Y10VDD_X70Y10VSS X70Y10VDDDM X70Y10VSS 0
I_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VDDDM 1 AC=0.006944444444444444
V_X70Y20VDD_X70Y20VSS X70Y20VDDDM X70Y20VSS 0
I_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VDDDM 1 AC=0.006944444444444444
V_X70Y30VDD_X70Y30VSS X70Y30VDDDM X70Y30VSS 0
I_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VDDDM 1 AC=0.006944444444444444
V_X70Y40VDD_X70Y40VSS X70Y40VDDDM X70Y40VSS 0
I_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VDDDM 1 AC=0.006944444444444444
V_X70Y50VDD_X70Y50VSS X70Y50VDDDM X70Y50VSS 0
I_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VDDDM 1 AC=0.006944444444444444
V_X70Y60VDD_X70Y60VSS X70Y60VDDDM X70Y60VSS 0
I_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VDDDM 1 AC=0.006944444444444444
V_X70Y70VDD_X70Y70VSS X70Y70VDDDM X70Y70VSS 0
I_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VDDDM 1 AC=0.006944444444444444
V_X70Y80VDD_X70Y80VSS X70Y80VDDDM X70Y80VSS 0
I_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VDDDM 1 AC=0.006944444444444444
V_X70Y90VDD_X70Y90VSS X70Y90VDDDM X70Y90VSS 0
I_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VDDDM 1 AC=0.006944444444444444
V_X70Y100VDD_X70Y100VSS X70Y100VDDDM X70Y100VSS 0
I_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VDDDM 1 AC=0.006944444444444444
V_X70Y110VDD_X70Y110VSS X70Y110VDDDM X70Y110VSS 0
I_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VDDDM 1 AC=0.006944444444444444
V_X80Y120VDD_X80Y120VSS X80Y120VDDDM X80Y120VSS 0
I_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VDDDM 1 AC=0.006944444444444444
V_X80Y10VDD_X80Y10VSS X80Y10VDDDM X80Y10VSS 0
I_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VDDDM 1 AC=0.006944444444444444
V_X80Y20VDD_X80Y20VSS X80Y20VDDDM X80Y20VSS 0
I_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VDDDM 1 AC=0.006944444444444444
V_X80Y30VDD_X80Y30VSS X80Y30VDDDM X80Y30VSS 0
I_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VDDDM 1 AC=0.006944444444444444
V_X80Y40VDD_X80Y40VSS X80Y40VDDDM X80Y40VSS 0
I_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VDDDM 1 AC=0.006944444444444444
V_X80Y50VDD_X80Y50VSS X80Y50VDDDM X80Y50VSS 0
I_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VDDDM 1 AC=0.006944444444444444
V_X80Y60VDD_X80Y60VSS X80Y60VDDDM X80Y60VSS 0
I_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VDDDM 1 AC=0.006944444444444444
V_X80Y70VDD_X80Y70VSS X80Y70VDDDM X80Y70VSS 0
I_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VDDDM 1 AC=0.006944444444444444
V_X80Y80VDD_X80Y80VSS X80Y80VDDDM X80Y80VSS 0
I_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VDDDM 1 AC=0.006944444444444444
V_X80Y90VDD_X80Y90VSS X80Y90VDDDM X80Y90VSS 0
I_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VDDDM 1 AC=0.006944444444444444
V_X80Y100VDD_X80Y100VSS X80Y100VDDDM X80Y100VSS 0
I_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VDDDM 1 AC=0.006944444444444444
V_X80Y110VDD_X80Y110VSS X80Y110VDDDM X80Y110VSS 0
I_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VDDDM 1 AC=0.006944444444444444
V_X90Y120VDD_X90Y120VSS X90Y120VDDDM X90Y120VSS 0
I_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VDDDM 1 AC=0.006944444444444444
V_X90Y10VDD_X90Y10VSS X90Y10VDDDM X90Y10VSS 0
I_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VDDDM 1 AC=0.006944444444444444
V_X90Y20VDD_X90Y20VSS X90Y20VDDDM X90Y20VSS 0
I_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VDDDM 1 AC=0.006944444444444444
V_X90Y30VDD_X90Y30VSS X90Y30VDDDM X90Y30VSS 0
I_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VDDDM 1 AC=0.006944444444444444
V_X90Y40VDD_X90Y40VSS X90Y40VDDDM X90Y40VSS 0
I_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VDDDM 1 AC=0.006944444444444444
V_X90Y50VDD_X90Y50VSS X90Y50VDDDM X90Y50VSS 0
I_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VDDDM 1 AC=0.006944444444444444
V_X90Y60VDD_X90Y60VSS X90Y60VDDDM X90Y60VSS 0
I_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VDDDM 1 AC=0.006944444444444444
V_X90Y70VDD_X90Y70VSS X90Y70VDDDM X90Y70VSS 0
I_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VDDDM 1 AC=0.006944444444444444
V_X90Y80VDD_X90Y80VSS X90Y80VDDDM X90Y80VSS 0
I_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VDDDM 1 AC=0.006944444444444444
V_X90Y90VDD_X90Y90VSS X90Y90VDDDM X90Y90VSS 0
I_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VDDDM 1 AC=0.006944444444444444
V_X90Y100VDD_X90Y100VSS X90Y100VDDDM X90Y100VSS 0
I_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VDDDM 1 AC=0.006944444444444444
V_X90Y110VDD_X90Y110VSS X90Y110VDDDM X90Y110VSS 0
I_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VDDDM 1 AC=0.006944444444444444
V_X100Y120VDD_X100Y120VSS X100Y120VDDDM X100Y120VSS 0
I_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VDDDM 1 AC=0.006944444444444444
V_X100Y10VDD_X100Y10VSS X100Y10VDDDM X100Y10VSS 0
I_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VDDDM 1 AC=0.006944444444444444
V_X100Y20VDD_X100Y20VSS X100Y20VDDDM X100Y20VSS 0
I_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VDDDM 1 AC=0.006944444444444444
V_X100Y30VDD_X100Y30VSS X100Y30VDDDM X100Y30VSS 0
I_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VDDDM 1 AC=0.006944444444444444
V_X100Y40VDD_X100Y40VSS X100Y40VDDDM X100Y40VSS 0
I_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VDDDM 1 AC=0.006944444444444444
V_X100Y50VDD_X100Y50VSS X100Y50VDDDM X100Y50VSS 0
I_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VDDDM 1 AC=0.006944444444444444
V_X100Y60VDD_X100Y60VSS X100Y60VDDDM X100Y60VSS 0
I_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VDDDM 1 AC=0.006944444444444444
V_X100Y70VDD_X100Y70VSS X100Y70VDDDM X100Y70VSS 0
I_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VDDDM 1 AC=0.006944444444444444
V_X100Y80VDD_X100Y80VSS X100Y80VDDDM X100Y80VSS 0
I_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VDDDM 1 AC=0.006944444444444444
V_X100Y90VDD_X100Y90VSS X100Y90VDDDM X100Y90VSS 0
I_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VDDDM 1 AC=0.006944444444444444
V_X100Y100VDD_X100Y100VSS X100Y100VDDDM X100Y100VSS 0
I_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VDDDM 1 AC=0.006944444444444444
V_X100Y110VDD_X100Y110VSS X100Y110VDDDM X100Y110VSS 0
I_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VDDDM 1 AC=0.006944444444444444
V_X110Y120VDD_X110Y120VSS X110Y120VDDDM X110Y120VSS 0
I_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VDDDM 1 AC=0.006944444444444444
V_X110Y10VDD_X110Y10VSS X110Y10VDDDM X110Y10VSS 0
I_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VDDDM 1 AC=0.006944444444444444
V_X110Y20VDD_X110Y20VSS X110Y20VDDDM X110Y20VSS 0
I_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VDDDM 1 AC=0.006944444444444444
V_X110Y30VDD_X110Y30VSS X110Y30VDDDM X110Y30VSS 0
I_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VDDDM 1 AC=0.006944444444444444
V_X110Y40VDD_X110Y40VSS X110Y40VDDDM X110Y40VSS 0
I_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VDDDM 1 AC=0.006944444444444444
V_X110Y50VDD_X110Y50VSS X110Y50VDDDM X110Y50VSS 0
I_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VDDDM 1 AC=0.006944444444444444
V_X110Y60VDD_X110Y60VSS X110Y60VDDDM X110Y60VSS 0
I_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VDDDM 1 AC=0.006944444444444444
V_X110Y70VDD_X110Y70VSS X110Y70VDDDM X110Y70VSS 0
I_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VDDDM 1 AC=0.006944444444444444
V_X110Y80VDD_X110Y80VSS X110Y80VDDDM X110Y80VSS 0
I_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VDDDM 1 AC=0.006944444444444444
V_X110Y90VDD_X110Y90VSS X110Y90VDDDM X110Y90VSS 0
I_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VDDDM 1 AC=0.006944444444444444
V_X110Y100VDD_X110Y100VSS X110Y100VDDDM X110Y100VSS 0
I_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VDDDM 1 AC=0.006944444444444444
V_X110Y110VDD_X110Y110VSS X110Y110VDDDM X110Y110VSS 0
Rbump_X10Y10VDD X10Y10VDD X10Y10VDDM 20mOhm
Lbump_X10Y10VDD X10Y10VDDM VDD2 0.036nH
Rbump_X10Y10VSS X10Y10VSS X10Y10VSSM 20mOhm
Lbump_X10Y10VSS X10Y10VSSM VSS2 0.036nH
Rbump_X10Y20VDD X10Y20VDD X10Y20VDDM 20mOhm
Lbump_X10Y20VDD X10Y20VDDM VDD2 0.036nH
Rbump_X10Y20VSS X10Y20VSS X10Y20VSSM 20mOhm
Lbump_X10Y20VSS X10Y20VSSM VSS2 0.036nH
Rbump_X10Y30VDD X10Y30VDD X10Y30VDDM 20mOhm
Lbump_X10Y30VDD X10Y30VDDM VDD2 0.036nH
Rbump_X10Y30VSS X10Y30VSS X10Y30VSSM 20mOhm
Lbump_X10Y30VSS X10Y30VSSM VSS2 0.036nH
Rbump_X10Y40VDD X10Y40VDD X10Y40VDDM 20mOhm
Lbump_X10Y40VDD X10Y40VDDM VDD2 0.036nH
Rbump_X10Y40VSS X10Y40VSS X10Y40VSSM 20mOhm
Lbump_X10Y40VSS X10Y40VSSM VSS2 0.036nH
Rbump_X10Y50VDD X10Y50VDD X10Y50VDDM 20mOhm
Lbump_X10Y50VDD X10Y50VDDM VDD2 0.036nH
Rbump_X10Y50VSS X10Y50VSS X10Y50VSSM 20mOhm
Lbump_X10Y50VSS X10Y50VSSM VSS2 0.036nH
Rbump_X10Y60VDD X10Y60VDD X10Y60VDDM 20mOhm
Lbump_X10Y60VDD X10Y60VDDM VDD2 0.036nH
Rbump_X10Y60VSS X10Y60VSS X10Y60VSSM 20mOhm
Lbump_X10Y60VSS X10Y60VSSM VSS2 0.036nH
Rbump_X10Y70VDD X10Y70VDD X10Y70VDDM 20mOhm
Lbump_X10Y70VDD X10Y70VDDM VDD2 0.036nH
Rbump_X10Y70VSS X10Y70VSS X10Y70VSSM 20mOhm
Lbump_X10Y70VSS X10Y70VSSM VSS2 0.036nH
Rbump_X10Y80VDD X10Y80VDD X10Y80VDDM 20mOhm
Lbump_X10Y80VDD X10Y80VDDM VDD2 0.036nH
Rbump_X10Y80VSS X10Y80VSS X10Y80VSSM 20mOhm
Lbump_X10Y80VSS X10Y80VSSM VSS2 0.036nH
Rbump_X10Y90VDD X10Y90VDD X10Y90VDDM 20mOhm
Lbump_X10Y90VDD X10Y90VDDM VDD2 0.036nH
Rbump_X10Y90VSS X10Y90VSS X10Y90VSSM 20mOhm
Lbump_X10Y90VSS X10Y90VSSM VSS2 0.036nH
Rbump_X10Y100VDD X10Y100VDD X10Y100VDDM 20mOhm
Lbump_X10Y100VDD X10Y100VDDM VDD2 0.036nH
Rbump_X10Y100VSS X10Y100VSS X10Y100VSSM 20mOhm
Lbump_X10Y100VSS X10Y100VSSM VSS2 0.036nH
Rbump_X10Y110VDD X10Y110VDD X10Y110VDDM 20mOhm
Lbump_X10Y110VDD X10Y110VDDM VDD2 0.036nH
Rbump_X10Y110VSS X10Y110VSS X10Y110VSSM 20mOhm
Lbump_X10Y110VSS X10Y110VSSM VSS2 0.036nH
Rbump_X10Y120VDD X10Y120VDD X10Y120VDDM 20mOhm
Lbump_X10Y120VDD X10Y120VDDM VDD2 0.036nH
Rbump_X10Y120VSS X10Y120VSS X10Y120VSSM 20mOhm
Lbump_X10Y120VSS X10Y120VSSM VSS2 0.036nH
Rbump_X20Y10VDD X20Y10VDD X20Y10VDDM 20mOhm
Lbump_X20Y10VDD X20Y10VDDM VDD2 0.036nH
Rbump_X20Y10VSS X20Y10VSS X20Y10VSSM 20mOhm
Lbump_X20Y10VSS X20Y10VSSM VSS2 0.036nH
Rbump_X20Y20VDD X20Y20VDD X20Y20VDDM 20mOhm
Lbump_X20Y20VDD X20Y20VDDM VDD2 0.036nH
Rbump_X20Y20VSS X20Y20VSS X20Y20VSSM 20mOhm
Lbump_X20Y20VSS X20Y20VSSM VSS2 0.036nH
Rbump_X20Y30VDD X20Y30VDD X20Y30VDDM 20mOhm
Lbump_X20Y30VDD X20Y30VDDM VDD2 0.036nH
Rbump_X20Y30VSS X20Y30VSS X20Y30VSSM 20mOhm
Lbump_X20Y30VSS X20Y30VSSM VSS2 0.036nH
Rbump_X20Y40VDD X20Y40VDD X20Y40VDDM 20mOhm
Lbump_X20Y40VDD X20Y40VDDM VDD2 0.036nH
Rbump_X20Y40VSS X20Y40VSS X20Y40VSSM 20mOhm
Lbump_X20Y40VSS X20Y40VSSM VSS2 0.036nH
Rbump_X20Y50VDD X20Y50VDD X20Y50VDDM 20mOhm
Lbump_X20Y50VDD X20Y50VDDM VDD2 0.036nH
Rbump_X20Y50VSS X20Y50VSS X20Y50VSSM 20mOhm
Lbump_X20Y50VSS X20Y50VSSM VSS2 0.036nH
Rbump_X20Y60VDD X20Y60VDD X20Y60VDDM 20mOhm
Lbump_X20Y60VDD X20Y60VDDM VDD2 0.036nH
Rbump_X20Y60VSS X20Y60VSS X20Y60VSSM 20mOhm
Lbump_X20Y60VSS X20Y60VSSM VSS2 0.036nH
Rbump_X20Y70VDD X20Y70VDD X20Y70VDDM 20mOhm
Lbump_X20Y70VDD X20Y70VDDM VDD2 0.036nH
Rbump_X20Y70VSS X20Y70VSS X20Y70VSSM 20mOhm
Lbump_X20Y70VSS X20Y70VSSM VSS2 0.036nH
Rbump_X20Y80VDD X20Y80VDD X20Y80VDDM 20mOhm
Lbump_X20Y80VDD X20Y80VDDM VDD2 0.036nH
Rbump_X20Y80VSS X20Y80VSS X20Y80VSSM 20mOhm
Lbump_X20Y80VSS X20Y80VSSM VSS2 0.036nH
Rbump_X20Y90VDD X20Y90VDD X20Y90VDDM 20mOhm
Lbump_X20Y90VDD X20Y90VDDM VDD2 0.036nH
Rbump_X20Y90VSS X20Y90VSS X20Y90VSSM 20mOhm
Lbump_X20Y90VSS X20Y90VSSM VSS2 0.036nH
Rbump_X20Y100VDD X20Y100VDD X20Y100VDDM 20mOhm
Lbump_X20Y100VDD X20Y100VDDM VDD2 0.036nH
Rbump_X20Y100VSS X20Y100VSS X20Y100VSSM 20mOhm
Lbump_X20Y100VSS X20Y100VSSM VSS2 0.036nH
Rbump_X20Y110VDD X20Y110VDD X20Y110VDDM 20mOhm
Lbump_X20Y110VDD X20Y110VDDM VDD2 0.036nH
Rbump_X20Y110VSS X20Y110VSS X20Y110VSSM 20mOhm
Lbump_X20Y110VSS X20Y110VSSM VSS2 0.036nH
Rbump_X20Y120VDD X20Y120VDD X20Y120VDDM 20mOhm
Lbump_X20Y120VDD X20Y120VDDM VDD2 0.036nH
Rbump_X20Y120VSS X20Y120VSS X20Y120VSSM 20mOhm
Lbump_X20Y120VSS X20Y120VSSM VSS2 0.036nH
Rbump_X30Y10VDD X30Y10VDD X30Y10VDDM 20mOhm
Lbump_X30Y10VDD X30Y10VDDM VDD2 0.036nH
Rbump_X30Y10VSS X30Y10VSS X30Y10VSSM 20mOhm
Lbump_X30Y10VSS X30Y10VSSM VSS2 0.036nH
Rbump_X30Y20VDD X30Y20VDD X30Y20VDDM 20mOhm
Lbump_X30Y20VDD X30Y20VDDM VDD2 0.036nH
Rbump_X30Y20VSS X30Y20VSS X30Y20VSSM 20mOhm
Lbump_X30Y20VSS X30Y20VSSM VSS2 0.036nH
Rbump_X30Y30VDD X30Y30VDD X30Y30VDDM 20mOhm
Lbump_X30Y30VDD X30Y30VDDM VDD2 0.036nH
Rbump_X30Y30VSS X30Y30VSS X30Y30VSSM 20mOhm
Lbump_X30Y30VSS X30Y30VSSM VSS2 0.036nH
Rbump_X30Y40VDD X30Y40VDD X30Y40VDDM 20mOhm
Lbump_X30Y40VDD X30Y40VDDM VDD2 0.036nH
Rbump_X30Y40VSS X30Y40VSS X30Y40VSSM 20mOhm
Lbump_X30Y40VSS X30Y40VSSM VSS2 0.036nH
Rbump_X30Y50VDD X30Y50VDD X30Y50VDDM 20mOhm
Lbump_X30Y50VDD X30Y50VDDM VDD2 0.036nH
Rbump_X30Y50VSS X30Y50VSS X30Y50VSSM 20mOhm
Lbump_X30Y50VSS X30Y50VSSM VSS2 0.036nH
Rbump_X30Y60VDD X30Y60VDD X30Y60VDDM 20mOhm
Lbump_X30Y60VDD X30Y60VDDM VDD2 0.036nH
Rbump_X30Y60VSS X30Y60VSS X30Y60VSSM 20mOhm
Lbump_X30Y60VSS X30Y60VSSM VSS2 0.036nH
Rbump_X30Y70VDD X30Y70VDD X30Y70VDDM 20mOhm
Lbump_X30Y70VDD X30Y70VDDM VDD2 0.036nH
Rbump_X30Y70VSS X30Y70VSS X30Y70VSSM 20mOhm
Lbump_X30Y70VSS X30Y70VSSM VSS2 0.036nH
Rbump_X30Y80VDD X30Y80VDD X30Y80VDDM 20mOhm
Lbump_X30Y80VDD X30Y80VDDM VDD2 0.036nH
Rbump_X30Y80VSS X30Y80VSS X30Y80VSSM 20mOhm
Lbump_X30Y80VSS X30Y80VSSM VSS2 0.036nH
Rbump_X30Y90VDD X30Y90VDD X30Y90VDDM 20mOhm
Lbump_X30Y90VDD X30Y90VDDM VDD2 0.036nH
Rbump_X30Y90VSS X30Y90VSS X30Y90VSSM 20mOhm
Lbump_X30Y90VSS X30Y90VSSM VSS2 0.036nH
Rbump_X30Y100VDD X30Y100VDD X30Y100VDDM 20mOhm
Lbump_X30Y100VDD X30Y100VDDM VDD2 0.036nH
Rbump_X30Y100VSS X30Y100VSS X30Y100VSSM 20mOhm
Lbump_X30Y100VSS X30Y100VSSM VSS2 0.036nH
Rbump_X30Y110VDD X30Y110VDD X30Y110VDDM 20mOhm
Lbump_X30Y110VDD X30Y110VDDM VDD2 0.036nH
Rbump_X30Y110VSS X30Y110VSS X30Y110VSSM 20mOhm
Lbump_X30Y110VSS X30Y110VSSM VSS2 0.036nH
Rbump_X30Y120VDD X30Y120VDD X30Y120VDDM 20mOhm
Lbump_X30Y120VDD X30Y120VDDM VDD2 0.036nH
Rbump_X30Y120VSS X30Y120VSS X30Y120VSSM 20mOhm
Lbump_X30Y120VSS X30Y120VSSM VSS2 0.036nH
Rbump_X40Y10VDD X40Y10VDD X40Y10VDDM 20mOhm
Lbump_X40Y10VDD X40Y10VDDM VDD2 0.036nH
Rbump_X40Y10VSS X40Y10VSS X40Y10VSSM 20mOhm
Lbump_X40Y10VSS X40Y10VSSM VSS2 0.036nH
Rbump_X40Y20VDD X40Y20VDD X40Y20VDDM 20mOhm
Lbump_X40Y20VDD X40Y20VDDM VDD2 0.036nH
Rbump_X40Y20VSS X40Y20VSS X40Y20VSSM 20mOhm
Lbump_X40Y20VSS X40Y20VSSM VSS2 0.036nH
Rbump_X40Y30VDD X40Y30VDD X40Y30VDDM 20mOhm
Lbump_X40Y30VDD X40Y30VDDM VDD2 0.036nH
Rbump_X40Y30VSS X40Y30VSS X40Y30VSSM 20mOhm
Lbump_X40Y30VSS X40Y30VSSM VSS2 0.036nH
Rbump_X40Y40VDD X40Y40VDD X40Y40VDDM 20mOhm
Lbump_X40Y40VDD X40Y40VDDM VDD2 0.036nH
Rbump_X40Y40VSS X40Y40VSS X40Y40VSSM 20mOhm
Lbump_X40Y40VSS X40Y40VSSM VSS2 0.036nH
Rbump_X40Y50VDD X40Y50VDD X40Y50VDDM 20mOhm
Lbump_X40Y50VDD X40Y50VDDM VDD2 0.036nH
Rbump_X40Y50VSS X40Y50VSS X40Y50VSSM 20mOhm
Lbump_X40Y50VSS X40Y50VSSM VSS2 0.036nH
Rbump_X40Y60VDD X40Y60VDD X40Y60VDDM 20mOhm
Lbump_X40Y60VDD X40Y60VDDM VDD2 0.036nH
Rbump_X40Y60VSS X40Y60VSS X40Y60VSSM 20mOhm
Lbump_X40Y60VSS X40Y60VSSM VSS2 0.036nH
Rbump_X40Y70VDD X40Y70VDD X40Y70VDDM 20mOhm
Lbump_X40Y70VDD X40Y70VDDM VDD2 0.036nH
Rbump_X40Y70VSS X40Y70VSS X40Y70VSSM 20mOhm
Lbump_X40Y70VSS X40Y70VSSM VSS2 0.036nH
Rbump_X40Y80VDD X40Y80VDD X40Y80VDDM 20mOhm
Lbump_X40Y80VDD X40Y80VDDM VDD2 0.036nH
Rbump_X40Y80VSS X40Y80VSS X40Y80VSSM 20mOhm
Lbump_X40Y80VSS X40Y80VSSM VSS2 0.036nH
Rbump_X40Y90VDD X40Y90VDD X40Y90VDDM 20mOhm
Lbump_X40Y90VDD X40Y90VDDM VDD2 0.036nH
Rbump_X40Y90VSS X40Y90VSS X40Y90VSSM 20mOhm
Lbump_X40Y90VSS X40Y90VSSM VSS2 0.036nH
Rbump_X40Y100VDD X40Y100VDD X40Y100VDDM 20mOhm
Lbump_X40Y100VDD X40Y100VDDM VDD2 0.036nH
Rbump_X40Y100VSS X40Y100VSS X40Y100VSSM 20mOhm
Lbump_X40Y100VSS X40Y100VSSM VSS2 0.036nH
Rbump_X40Y110VDD X40Y110VDD X40Y110VDDM 20mOhm
Lbump_X40Y110VDD X40Y110VDDM VDD2 0.036nH
Rbump_X40Y110VSS X40Y110VSS X40Y110VSSM 20mOhm
Lbump_X40Y110VSS X40Y110VSSM VSS2 0.036nH
Rbump_X40Y120VDD X40Y120VDD X40Y120VDDM 20mOhm
Lbump_X40Y120VDD X40Y120VDDM VDD2 0.036nH
Rbump_X40Y120VSS X40Y120VSS X40Y120VSSM 20mOhm
Lbump_X40Y120VSS X40Y120VSSM VSS2 0.036nH
Rbump_X50Y10VDD X50Y10VDD X50Y10VDDM 20mOhm
Lbump_X50Y10VDD X50Y10VDDM VDD2 0.036nH
Rbump_X50Y10VSS X50Y10VSS X50Y10VSSM 20mOhm
Lbump_X50Y10VSS X50Y10VSSM VSS2 0.036nH
Rbump_X50Y20VDD X50Y20VDD X50Y20VDDM 20mOhm
Lbump_X50Y20VDD X50Y20VDDM VDD2 0.036nH
Rbump_X50Y20VSS X50Y20VSS X50Y20VSSM 20mOhm
Lbump_X50Y20VSS X50Y20VSSM VSS2 0.036nH
Rbump_X50Y30VDD X50Y30VDD X50Y30VDDM 20mOhm
Lbump_X50Y30VDD X50Y30VDDM VDD2 0.036nH
Rbump_X50Y30VSS X50Y30VSS X50Y30VSSM 20mOhm
Lbump_X50Y30VSS X50Y30VSSM VSS2 0.036nH
Rbump_X50Y40VDD X50Y40VDD X50Y40VDDM 20mOhm
Lbump_X50Y40VDD X50Y40VDDM VDD2 0.036nH
Rbump_X50Y40VSS X50Y40VSS X50Y40VSSM 20mOhm
Lbump_X50Y40VSS X50Y40VSSM VSS2 0.036nH
Rbump_X50Y50VDD X50Y50VDD X50Y50VDDM 20mOhm
Lbump_X50Y50VDD X50Y50VDDM VDD2 0.036nH
Rbump_X50Y50VSS X50Y50VSS X50Y50VSSM 20mOhm
Lbump_X50Y50VSS X50Y50VSSM VSS2 0.036nH
Rbump_X50Y60VDD X50Y60VDD X50Y60VDDM 20mOhm
Lbump_X50Y60VDD X50Y60VDDM VDD2 0.036nH
Rbump_X50Y60VSS X50Y60VSS X50Y60VSSM 20mOhm
Lbump_X50Y60VSS X50Y60VSSM VSS2 0.036nH
Rbump_X50Y70VDD X50Y70VDD X50Y70VDDM 20mOhm
Lbump_X50Y70VDD X50Y70VDDM VDD2 0.036nH
Rbump_X50Y70VSS X50Y70VSS X50Y70VSSM 20mOhm
Lbump_X50Y70VSS X50Y70VSSM VSS2 0.036nH
Rbump_X50Y80VDD X50Y80VDD X50Y80VDDM 20mOhm
Lbump_X50Y80VDD X50Y80VDDM VDD2 0.036nH
Rbump_X50Y80VSS X50Y80VSS X50Y80VSSM 20mOhm
Lbump_X50Y80VSS X50Y80VSSM VSS2 0.036nH
Rbump_X50Y90VDD X50Y90VDD X50Y90VDDM 20mOhm
Lbump_X50Y90VDD X50Y90VDDM VDD2 0.036nH
Rbump_X50Y90VSS X50Y90VSS X50Y90VSSM 20mOhm
Lbump_X50Y90VSS X50Y90VSSM VSS2 0.036nH
Rbump_X50Y100VDD X50Y100VDD X50Y100VDDM 20mOhm
Lbump_X50Y100VDD X50Y100VDDM VDD2 0.036nH
Rbump_X50Y100VSS X50Y100VSS X50Y100VSSM 20mOhm
Lbump_X50Y100VSS X50Y100VSSM VSS2 0.036nH
Rbump_X50Y110VDD X50Y110VDD X50Y110VDDM 20mOhm
Lbump_X50Y110VDD X50Y110VDDM VDD2 0.036nH
Rbump_X50Y110VSS X50Y110VSS X50Y110VSSM 20mOhm
Lbump_X50Y110VSS X50Y110VSSM VSS2 0.036nH
Rbump_X50Y120VDD X50Y120VDD X50Y120VDDM 20mOhm
Lbump_X50Y120VDD X50Y120VDDM VDD2 0.036nH
Rbump_X50Y120VSS X50Y120VSS X50Y120VSSM 20mOhm
Lbump_X50Y120VSS X50Y120VSSM VSS2 0.036nH
Rbump_X60Y10VDD X60Y10VDD X60Y10VDDM 20mOhm
Lbump_X60Y10VDD X60Y10VDDM VDD2 0.036nH
Rbump_X60Y10VSS X60Y10VSS X60Y10VSSM 20mOhm
Lbump_X60Y10VSS X60Y10VSSM VSS2 0.036nH
Rbump_X60Y20VDD X60Y20VDD X60Y20VDDM 20mOhm
Lbump_X60Y20VDD X60Y20VDDM VDD2 0.036nH
Rbump_X60Y20VSS X60Y20VSS X60Y20VSSM 20mOhm
Lbump_X60Y20VSS X60Y20VSSM VSS2 0.036nH
Rbump_X60Y30VDD X60Y30VDD X60Y30VDDM 20mOhm
Lbump_X60Y30VDD X60Y30VDDM VDD2 0.036nH
Rbump_X60Y30VSS X60Y30VSS X60Y30VSSM 20mOhm
Lbump_X60Y30VSS X60Y30VSSM VSS2 0.036nH
Rbump_X60Y40VDD X60Y40VDD X60Y40VDDM 20mOhm
Lbump_X60Y40VDD X60Y40VDDM VDD2 0.036nH
Rbump_X60Y40VSS X60Y40VSS X60Y40VSSM 20mOhm
Lbump_X60Y40VSS X60Y40VSSM VSS2 0.036nH
Rbump_X60Y50VDD X60Y50VDD X60Y50VDDM 20mOhm
Lbump_X60Y50VDD X60Y50VDDM VDD2 0.036nH
Rbump_X60Y50VSS X60Y50VSS X60Y50VSSM 20mOhm
Lbump_X60Y50VSS X60Y50VSSM VSS2 0.036nH
Rbump_X60Y60VDD X60Y60VDD X60Y60VDDM 20mOhm
Lbump_X60Y60VDD X60Y60VDDM VDD2 0.036nH
Rbump_X60Y60VSS X60Y60VSS X60Y60VSSM 20mOhm
Lbump_X60Y60VSS X60Y60VSSM VSS2 0.036nH
Rbump_X60Y70VDD X60Y70VDD X60Y70VDDM 20mOhm
Lbump_X60Y70VDD X60Y70VDDM VDD2 0.036nH
Rbump_X60Y70VSS X60Y70VSS X60Y70VSSM 20mOhm
Lbump_X60Y70VSS X60Y70VSSM VSS2 0.036nH
Rbump_X60Y80VDD X60Y80VDD X60Y80VDDM 20mOhm
Lbump_X60Y80VDD X60Y80VDDM VDD2 0.036nH
Rbump_X60Y80VSS X60Y80VSS X60Y80VSSM 20mOhm
Lbump_X60Y80VSS X60Y80VSSM VSS2 0.036nH
Rbump_X60Y90VDD X60Y90VDD X60Y90VDDM 20mOhm
Lbump_X60Y90VDD X60Y90VDDM VDD2 0.036nH
Rbump_X60Y90VSS X60Y90VSS X60Y90VSSM 20mOhm
Lbump_X60Y90VSS X60Y90VSSM VSS2 0.036nH
Rbump_X60Y100VDD X60Y100VDD X60Y100VDDM 20mOhm
Lbump_X60Y100VDD X60Y100VDDM VDD2 0.036nH
Rbump_X60Y100VSS X60Y100VSS X60Y100VSSM 20mOhm
Lbump_X60Y100VSS X60Y100VSSM VSS2 0.036nH
Rbump_X60Y110VDD X60Y110VDD X60Y110VDDM 20mOhm
Lbump_X60Y110VDD X60Y110VDDM VDD2 0.036nH
Rbump_X60Y110VSS X60Y110VSS X60Y110VSSM 20mOhm
Lbump_X60Y110VSS X60Y110VSSM VSS2 0.036nH
Rbump_X60Y120VDD X60Y120VDD X60Y120VDDM 20mOhm
Lbump_X60Y120VDD X60Y120VDDM VDD2 0.036nH
Rbump_X60Y120VSS X60Y120VSS X60Y120VSSM 20mOhm
Lbump_X60Y120VSS X60Y120VSSM VSS2 0.036nH
Rbump_X70Y10VDD X70Y10VDD X70Y10VDDM 20mOhm
Lbump_X70Y10VDD X70Y10VDDM VDD2 0.036nH
Rbump_X70Y10VSS X70Y10VSS X70Y10VSSM 20mOhm
Lbump_X70Y10VSS X70Y10VSSM VSS2 0.036nH
Rbump_X70Y20VDD X70Y20VDD X70Y20VDDM 20mOhm
Lbump_X70Y20VDD X70Y20VDDM VDD2 0.036nH
Rbump_X70Y20VSS X70Y20VSS X70Y20VSSM 20mOhm
Lbump_X70Y20VSS X70Y20VSSM VSS2 0.036nH
Rbump_X70Y30VDD X70Y30VDD X70Y30VDDM 20mOhm
Lbump_X70Y30VDD X70Y30VDDM VDD2 0.036nH
Rbump_X70Y30VSS X70Y30VSS X70Y30VSSM 20mOhm
Lbump_X70Y30VSS X70Y30VSSM VSS2 0.036nH
Rbump_X70Y40VDD X70Y40VDD X70Y40VDDM 20mOhm
Lbump_X70Y40VDD X70Y40VDDM VDD2 0.036nH
Rbump_X70Y40VSS X70Y40VSS X70Y40VSSM 20mOhm
Lbump_X70Y40VSS X70Y40VSSM VSS2 0.036nH
Rbump_X70Y50VDD X70Y50VDD X70Y50VDDM 20mOhm
Lbump_X70Y50VDD X70Y50VDDM VDD2 0.036nH
Rbump_X70Y50VSS X70Y50VSS X70Y50VSSM 20mOhm
Lbump_X70Y50VSS X70Y50VSSM VSS2 0.036nH
Rbump_X70Y60VDD X70Y60VDD X70Y60VDDM 20mOhm
Lbump_X70Y60VDD X70Y60VDDM VDD2 0.036nH
Rbump_X70Y60VSS X70Y60VSS X70Y60VSSM 20mOhm
Lbump_X70Y60VSS X70Y60VSSM VSS2 0.036nH
Rbump_X70Y70VDD X70Y70VDD X70Y70VDDM 20mOhm
Lbump_X70Y70VDD X70Y70VDDM VDD2 0.036nH
Rbump_X70Y70VSS X70Y70VSS X70Y70VSSM 20mOhm
Lbump_X70Y70VSS X70Y70VSSM VSS2 0.036nH
Rbump_X70Y80VDD X70Y80VDD X70Y80VDDM 20mOhm
Lbump_X70Y80VDD X70Y80VDDM VDD2 0.036nH
Rbump_X70Y80VSS X70Y80VSS X70Y80VSSM 20mOhm
Lbump_X70Y80VSS X70Y80VSSM VSS2 0.036nH
Rbump_X70Y90VDD X70Y90VDD X70Y90VDDM 20mOhm
Lbump_X70Y90VDD X70Y90VDDM VDD2 0.036nH
Rbump_X70Y90VSS X70Y90VSS X70Y90VSSM 20mOhm
Lbump_X70Y90VSS X70Y90VSSM VSS2 0.036nH
Rbump_X70Y100VDD X70Y100VDD X70Y100VDDM 20mOhm
Lbump_X70Y100VDD X70Y100VDDM VDD2 0.036nH
Rbump_X70Y100VSS X70Y100VSS X70Y100VSSM 20mOhm
Lbump_X70Y100VSS X70Y100VSSM VSS2 0.036nH
Rbump_X70Y110VDD X70Y110VDD X70Y110VDDM 20mOhm
Lbump_X70Y110VDD X70Y110VDDM VDD2 0.036nH
Rbump_X70Y110VSS X70Y110VSS X70Y110VSSM 20mOhm
Lbump_X70Y110VSS X70Y110VSSM VSS2 0.036nH
Rbump_X70Y120VDD X70Y120VDD X70Y120VDDM 20mOhm
Lbump_X70Y120VDD X70Y120VDDM VDD2 0.036nH
Rbump_X70Y120VSS X70Y120VSS X70Y120VSSM 20mOhm
Lbump_X70Y120VSS X70Y120VSSM VSS2 0.036nH
Rbump_X80Y10VDD X80Y10VDD X80Y10VDDM 20mOhm
Lbump_X80Y10VDD X80Y10VDDM VDD2 0.036nH
Rbump_X80Y10VSS X80Y10VSS X80Y10VSSM 20mOhm
Lbump_X80Y10VSS X80Y10VSSM VSS2 0.036nH
Rbump_X80Y20VDD X80Y20VDD X80Y20VDDM 20mOhm
Lbump_X80Y20VDD X80Y20VDDM VDD2 0.036nH
Rbump_X80Y20VSS X80Y20VSS X80Y20VSSM 20mOhm
Lbump_X80Y20VSS X80Y20VSSM VSS2 0.036nH
Rbump_X80Y30VDD X80Y30VDD X80Y30VDDM 20mOhm
Lbump_X80Y30VDD X80Y30VDDM VDD2 0.036nH
Rbump_X80Y30VSS X80Y30VSS X80Y30VSSM 20mOhm
Lbump_X80Y30VSS X80Y30VSSM VSS2 0.036nH
Rbump_X80Y40VDD X80Y40VDD X80Y40VDDM 20mOhm
Lbump_X80Y40VDD X80Y40VDDM VDD2 0.036nH
Rbump_X80Y40VSS X80Y40VSS X80Y40VSSM 20mOhm
Lbump_X80Y40VSS X80Y40VSSM VSS2 0.036nH
Rbump_X80Y50VDD X80Y50VDD X80Y50VDDM 20mOhm
Lbump_X80Y50VDD X80Y50VDDM VDD2 0.036nH
Rbump_X80Y50VSS X80Y50VSS X80Y50VSSM 20mOhm
Lbump_X80Y50VSS X80Y50VSSM VSS2 0.036nH
Rbump_X80Y60VDD X80Y60VDD X80Y60VDDM 20mOhm
Lbump_X80Y60VDD X80Y60VDDM VDD2 0.036nH
Rbump_X80Y60VSS X80Y60VSS X80Y60VSSM 20mOhm
Lbump_X80Y60VSS X80Y60VSSM VSS2 0.036nH
Rbump_X80Y70VDD X80Y70VDD X80Y70VDDM 20mOhm
Lbump_X80Y70VDD X80Y70VDDM VDD2 0.036nH
Rbump_X80Y70VSS X80Y70VSS X80Y70VSSM 20mOhm
Lbump_X80Y70VSS X80Y70VSSM VSS2 0.036nH
Rbump_X80Y80VDD X80Y80VDD X80Y80VDDM 20mOhm
Lbump_X80Y80VDD X80Y80VDDM VDD2 0.036nH
Rbump_X80Y80VSS X80Y80VSS X80Y80VSSM 20mOhm
Lbump_X80Y80VSS X80Y80VSSM VSS2 0.036nH
Rbump_X80Y90VDD X80Y90VDD X80Y90VDDM 20mOhm
Lbump_X80Y90VDD X80Y90VDDM VDD2 0.036nH
Rbump_X80Y90VSS X80Y90VSS X80Y90VSSM 20mOhm
Lbump_X80Y90VSS X80Y90VSSM VSS2 0.036nH
Rbump_X80Y100VDD X80Y100VDD X80Y100VDDM 20mOhm
Lbump_X80Y100VDD X80Y100VDDM VDD2 0.036nH
Rbump_X80Y100VSS X80Y100VSS X80Y100VSSM 20mOhm
Lbump_X80Y100VSS X80Y100VSSM VSS2 0.036nH
Rbump_X80Y110VDD X80Y110VDD X80Y110VDDM 20mOhm
Lbump_X80Y110VDD X80Y110VDDM VDD2 0.036nH
Rbump_X80Y110VSS X80Y110VSS X80Y110VSSM 20mOhm
Lbump_X80Y110VSS X80Y110VSSM VSS2 0.036nH
Rbump_X80Y120VDD X80Y120VDD X80Y120VDDM 20mOhm
Lbump_X80Y120VDD X80Y120VDDM VDD2 0.036nH
Rbump_X80Y120VSS X80Y120VSS X80Y120VSSM 20mOhm
Lbump_X80Y120VSS X80Y120VSSM VSS2 0.036nH
Rbump_X90Y10VDD X90Y10VDD X90Y10VDDM 20mOhm
Lbump_X90Y10VDD X90Y10VDDM VDD2 0.036nH
Rbump_X90Y10VSS X90Y10VSS X90Y10VSSM 20mOhm
Lbump_X90Y10VSS X90Y10VSSM VSS2 0.036nH
Rbump_X90Y20VDD X90Y20VDD X90Y20VDDM 20mOhm
Lbump_X90Y20VDD X90Y20VDDM VDD2 0.036nH
Rbump_X90Y20VSS X90Y20VSS X90Y20VSSM 20mOhm
Lbump_X90Y20VSS X90Y20VSSM VSS2 0.036nH
Rbump_X90Y30VDD X90Y30VDD X90Y30VDDM 20mOhm
Lbump_X90Y30VDD X90Y30VDDM VDD2 0.036nH
Rbump_X90Y30VSS X90Y30VSS X90Y30VSSM 20mOhm
Lbump_X90Y30VSS X90Y30VSSM VSS2 0.036nH
Rbump_X90Y40VDD X90Y40VDD X90Y40VDDM 20mOhm
Lbump_X90Y40VDD X90Y40VDDM VDD2 0.036nH
Rbump_X90Y40VSS X90Y40VSS X90Y40VSSM 20mOhm
Lbump_X90Y40VSS X90Y40VSSM VSS2 0.036nH
Rbump_X90Y50VDD X90Y50VDD X90Y50VDDM 20mOhm
Lbump_X90Y50VDD X90Y50VDDM VDD2 0.036nH
Rbump_X90Y50VSS X90Y50VSS X90Y50VSSM 20mOhm
Lbump_X90Y50VSS X90Y50VSSM VSS2 0.036nH
Rbump_X90Y60VDD X90Y60VDD X90Y60VDDM 20mOhm
Lbump_X90Y60VDD X90Y60VDDM VDD2 0.036nH
Rbump_X90Y60VSS X90Y60VSS X90Y60VSSM 20mOhm
Lbump_X90Y60VSS X90Y60VSSM VSS2 0.036nH
Rbump_X90Y70VDD X90Y70VDD X90Y70VDDM 20mOhm
Lbump_X90Y70VDD X90Y70VDDM VDD2 0.036nH
Rbump_X90Y70VSS X90Y70VSS X90Y70VSSM 20mOhm
Lbump_X90Y70VSS X90Y70VSSM VSS2 0.036nH
Rbump_X90Y80VDD X90Y80VDD X90Y80VDDM 20mOhm
Lbump_X90Y80VDD X90Y80VDDM VDD2 0.036nH
Rbump_X90Y80VSS X90Y80VSS X90Y80VSSM 20mOhm
Lbump_X90Y80VSS X90Y80VSSM VSS2 0.036nH
Rbump_X90Y90VDD X90Y90VDD X90Y90VDDM 20mOhm
Lbump_X90Y90VDD X90Y90VDDM VDD2 0.036nH
Rbump_X90Y90VSS X90Y90VSS X90Y90VSSM 20mOhm
Lbump_X90Y90VSS X90Y90VSSM VSS2 0.036nH
Rbump_X90Y100VDD X90Y100VDD X90Y100VDDM 20mOhm
Lbump_X90Y100VDD X90Y100VDDM VDD2 0.036nH
Rbump_X90Y100VSS X90Y100VSS X90Y100VSSM 20mOhm
Lbump_X90Y100VSS X90Y100VSSM VSS2 0.036nH
Rbump_X90Y110VDD X90Y110VDD X90Y110VDDM 20mOhm
Lbump_X90Y110VDD X90Y110VDDM VDD2 0.036nH
Rbump_X90Y110VSS X90Y110VSS X90Y110VSSM 20mOhm
Lbump_X90Y110VSS X90Y110VSSM VSS2 0.036nH
Rbump_X90Y120VDD X90Y120VDD X90Y120VDDM 20mOhm
Lbump_X90Y120VDD X90Y120VDDM VDD2 0.036nH
Rbump_X90Y120VSS X90Y120VSS X90Y120VSSM 20mOhm
Lbump_X90Y120VSS X90Y120VSSM VSS2 0.036nH
Rbump_X100Y10VDD X100Y10VDD X100Y10VDDM 20mOhm
Lbump_X100Y10VDD X100Y10VDDM VDD2 0.036nH
Rbump_X100Y10VSS X100Y10VSS X100Y10VSSM 20mOhm
Lbump_X100Y10VSS X100Y10VSSM VSS2 0.036nH
Rbump_X100Y20VDD X100Y20VDD X100Y20VDDM 20mOhm
Lbump_X100Y20VDD X100Y20VDDM VDD2 0.036nH
Rbump_X100Y20VSS X100Y20VSS X100Y20VSSM 20mOhm
Lbump_X100Y20VSS X100Y20VSSM VSS2 0.036nH
Rbump_X100Y30VDD X100Y30VDD X100Y30VDDM 20mOhm
Lbump_X100Y30VDD X100Y30VDDM VDD2 0.036nH
Rbump_X100Y30VSS X100Y30VSS X100Y30VSSM 20mOhm
Lbump_X100Y30VSS X100Y30VSSM VSS2 0.036nH
Rbump_X100Y40VDD X100Y40VDD X100Y40VDDM 20mOhm
Lbump_X100Y40VDD X100Y40VDDM VDD2 0.036nH
Rbump_X100Y40VSS X100Y40VSS X100Y40VSSM 20mOhm
Lbump_X100Y40VSS X100Y40VSSM VSS2 0.036nH
Rbump_X100Y50VDD X100Y50VDD X100Y50VDDM 20mOhm
Lbump_X100Y50VDD X100Y50VDDM VDD2 0.036nH
Rbump_X100Y50VSS X100Y50VSS X100Y50VSSM 20mOhm
Lbump_X100Y50VSS X100Y50VSSM VSS2 0.036nH
Rbump_X100Y60VDD X100Y60VDD X100Y60VDDM 20mOhm
Lbump_X100Y60VDD X100Y60VDDM VDD2 0.036nH
Rbump_X100Y60VSS X100Y60VSS X100Y60VSSM 20mOhm
Lbump_X100Y60VSS X100Y60VSSM VSS2 0.036nH
Rbump_X100Y70VDD X100Y70VDD X100Y70VDDM 20mOhm
Lbump_X100Y70VDD X100Y70VDDM VDD2 0.036nH
Rbump_X100Y70VSS X100Y70VSS X100Y70VSSM 20mOhm
Lbump_X100Y70VSS X100Y70VSSM VSS2 0.036nH
Rbump_X100Y80VDD X100Y80VDD X100Y80VDDM 20mOhm
Lbump_X100Y80VDD X100Y80VDDM VDD2 0.036nH
Rbump_X100Y80VSS X100Y80VSS X100Y80VSSM 20mOhm
Lbump_X100Y80VSS X100Y80VSSM VSS2 0.036nH
Rbump_X100Y90VDD X100Y90VDD X100Y90VDDM 20mOhm
Lbump_X100Y90VDD X100Y90VDDM VDD2 0.036nH
Rbump_X100Y90VSS X100Y90VSS X100Y90VSSM 20mOhm
Lbump_X100Y90VSS X100Y90VSSM VSS2 0.036nH
Rbump_X100Y100VDD X100Y100VDD X100Y100VDDM 20mOhm
Lbump_X100Y100VDD X100Y100VDDM VDD2 0.036nH
Rbump_X100Y100VSS X100Y100VSS X100Y100VSSM 20mOhm
Lbump_X100Y100VSS X100Y100VSSM VSS2 0.036nH
Rbump_X100Y110VDD X100Y110VDD X100Y110VDDM 20mOhm
Lbump_X100Y110VDD X100Y110VDDM VDD2 0.036nH
Rbump_X100Y110VSS X100Y110VSS X100Y110VSSM 20mOhm
Lbump_X100Y110VSS X100Y110VSSM VSS2 0.036nH
Rbump_X100Y120VDD X100Y120VDD X100Y120VDDM 20mOhm
Lbump_X100Y120VDD X100Y120VDDM VDD2 0.036nH
Rbump_X100Y120VSS X100Y120VSS X100Y120VSSM 20mOhm
Lbump_X100Y120VSS X100Y120VSSM VSS2 0.036nH
Rbump_X110Y10VDD X110Y10VDD X110Y10VDDM 20mOhm
Lbump_X110Y10VDD X110Y10VDDM VDD2 0.036nH
Rbump_X110Y10VSS X110Y10VSS X110Y10VSSM 20mOhm
Lbump_X110Y10VSS X110Y10VSSM VSS2 0.036nH
Rbump_X110Y20VDD X110Y20VDD X110Y20VDDM 20mOhm
Lbump_X110Y20VDD X110Y20VDDM VDD2 0.036nH
Rbump_X110Y20VSS X110Y20VSS X110Y20VSSM 20mOhm
Lbump_X110Y20VSS X110Y20VSSM VSS2 0.036nH
Rbump_X110Y30VDD X110Y30VDD X110Y30VDDM 20mOhm
Lbump_X110Y30VDD X110Y30VDDM VDD2 0.036nH
Rbump_X110Y30VSS X110Y30VSS X110Y30VSSM 20mOhm
Lbump_X110Y30VSS X110Y30VSSM VSS2 0.036nH
Rbump_X110Y40VDD X110Y40VDD X110Y40VDDM 20mOhm
Lbump_X110Y40VDD X110Y40VDDM VDD2 0.036nH
Rbump_X110Y40VSS X110Y40VSS X110Y40VSSM 20mOhm
Lbump_X110Y40VSS X110Y40VSSM VSS2 0.036nH
Rbump_X110Y50VDD X110Y50VDD X110Y50VDDM 20mOhm
Lbump_X110Y50VDD X110Y50VDDM VDD2 0.036nH
Rbump_X110Y50VSS X110Y50VSS X110Y50VSSM 20mOhm
Lbump_X110Y50VSS X110Y50VSSM VSS2 0.036nH
Rbump_X110Y60VDD X110Y60VDD X110Y60VDDM 20mOhm
Lbump_X110Y60VDD X110Y60VDDM VDD2 0.036nH
Rbump_X110Y60VSS X110Y60VSS X110Y60VSSM 20mOhm
Lbump_X110Y60VSS X110Y60VSSM VSS2 0.036nH
Rbump_X110Y70VDD X110Y70VDD X110Y70VDDM 20mOhm
Lbump_X110Y70VDD X110Y70VDDM VDD2 0.036nH
Rbump_X110Y70VSS X110Y70VSS X110Y70VSSM 20mOhm
Lbump_X110Y70VSS X110Y70VSSM VSS2 0.036nH
Rbump_X110Y80VDD X110Y80VDD X110Y80VDDM 20mOhm
Lbump_X110Y80VDD X110Y80VDDM VDD2 0.036nH
Rbump_X110Y80VSS X110Y80VSS X110Y80VSSM 20mOhm
Lbump_X110Y80VSS X110Y80VSSM VSS2 0.036nH
Rbump_X110Y90VDD X110Y90VDD X110Y90VDDM 20mOhm
Lbump_X110Y90VDD X110Y90VDDM VDD2 0.036nH
Rbump_X110Y90VSS X110Y90VSS X110Y90VSSM 20mOhm
Lbump_X110Y90VSS X110Y90VSSM VSS2 0.036nH
Rbump_X110Y100VDD X110Y100VDD X110Y100VDDM 20mOhm
Lbump_X110Y100VDD X110Y100VDDM VDD2 0.036nH
Rbump_X110Y100VSS X110Y100VSS X110Y100VSSM 20mOhm
Lbump_X110Y100VSS X110Y100VSSM VSS2 0.036nH
Rbump_X110Y110VDD X110Y110VDD X110Y110VDDM 20mOhm
Lbump_X110Y110VDD X110Y110VDDM VDD2 0.036nH
Rbump_X110Y110VSS X110Y110VSS X110Y110VSSM 20mOhm
Lbump_X110Y110VSS X110Y110VSSM VSS2 0.036nH
Rbump_X110Y120VDD X110Y120VDD X110Y120VDDM 20mOhm
Lbump_X110Y120VDD X110Y120VDDM VDD2 0.036nH
Rbump_X110Y120VSS X110Y120VSS X110Y120VSSM 20mOhm
Lbump_X110Y120VSS X110Y120VSSM VSS2 0.036nH
Rbump_X120Y10VDD X120Y10VDD X120Y10VDDM 20mOhm
Lbump_X120Y10VDD X120Y10VDDM VDD2 0.036nH
Rbump_X120Y10VSS X120Y10VSS X120Y10VSSM 20mOhm
Lbump_X120Y10VSS X120Y10VSSM VSS2 0.036nH
Rbump_X120Y20VDD X120Y20VDD X120Y20VDDM 20mOhm
Lbump_X120Y20VDD X120Y20VDDM VDD2 0.036nH
Rbump_X120Y20VSS X120Y20VSS X120Y20VSSM 20mOhm
Lbump_X120Y20VSS X120Y20VSSM VSS2 0.036nH
Rbump_X120Y30VDD X120Y30VDD X120Y30VDDM 20mOhm
Lbump_X120Y30VDD X120Y30VDDM VDD2 0.036nH
Rbump_X120Y30VSS X120Y30VSS X120Y30VSSM 20mOhm
Lbump_X120Y30VSS X120Y30VSSM VSS2 0.036nH
Rbump_X120Y40VDD X120Y40VDD X120Y40VDDM 20mOhm
Lbump_X120Y40VDD X120Y40VDDM VDD2 0.036nH
Rbump_X120Y40VSS X120Y40VSS X120Y40VSSM 20mOhm
Lbump_X120Y40VSS X120Y40VSSM VSS2 0.036nH
Rbump_X120Y50VDD X120Y50VDD X120Y50VDDM 20mOhm
Lbump_X120Y50VDD X120Y50VDDM VDD2 0.036nH
Rbump_X120Y50VSS X120Y50VSS X120Y50VSSM 20mOhm
Lbump_X120Y50VSS X120Y50VSSM VSS2 0.036nH
Rbump_X120Y60VDD X120Y60VDD X120Y60VDDM 20mOhm
Lbump_X120Y60VDD X120Y60VDDM VDD2 0.036nH
Rbump_X120Y60VSS X120Y60VSS X120Y60VSSM 20mOhm
Lbump_X120Y60VSS X120Y60VSSM VSS2 0.036nH
Rbump_X120Y70VDD X120Y70VDD X120Y70VDDM 20mOhm
Lbump_X120Y70VDD X120Y70VDDM VDD2 0.036nH
Rbump_X120Y70VSS X120Y70VSS X120Y70VSSM 20mOhm
Lbump_X120Y70VSS X120Y70VSSM VSS2 0.036nH
Rbump_X120Y80VDD X120Y80VDD X120Y80VDDM 20mOhm
Lbump_X120Y80VDD X120Y80VDDM VDD2 0.036nH
Rbump_X120Y80VSS X120Y80VSS X120Y80VSSM 20mOhm
Lbump_X120Y80VSS X120Y80VSSM VSS2 0.036nH
Rbump_X120Y90VDD X120Y90VDD X120Y90VDDM 20mOhm
Lbump_X120Y90VDD X120Y90VDDM VDD2 0.036nH
Rbump_X120Y90VSS X120Y90VSS X120Y90VSSM 20mOhm
Lbump_X120Y90VSS X120Y90VSSM VSS2 0.036nH
Rbump_X120Y100VDD X120Y100VDD X120Y100VDDM 20mOhm
Lbump_X120Y100VDD X120Y100VDDM VDD2 0.036nH
Rbump_X120Y100VSS X120Y100VSS X120Y100VSSM 20mOhm
Lbump_X120Y100VSS X120Y100VSSM VSS2 0.036nH
Rbump_X120Y110VDD X120Y110VDD X120Y110VDDM 20mOhm
Lbump_X120Y110VDD X120Y110VDDM VDD2 0.036nH
Rbump_X120Y110VSS X120Y110VSS X120Y110VSSM 20mOhm
Lbump_X120Y110VSS X120Y110VSSM VSS2 0.036nH
Rbump_X120Y120VDD X120Y120VDD X120Y120VDDM 20mOhm
Lbump_X120Y120VDD X120Y120VDDM VDD2 0.036nH
Rbump_X120Y120VSS X120Y120VSS X120Y120VSSM 20mOhm
Lbump_X120Y120VSS X120Y120VSSM VSS2 0.036nH
RsVDD VDD VDDMS 0.55mOhm
LsVDD VDDMS VDD2 0.06nH
RsVSS VSS VSSMS 0.55mOhm
LsVSS VSSMS VSS2 0.06nH
Rp VDD2 VDD2M 0.1mOhm
Lp VSS2 VSS2M 0.0028nH
Cp VDD2M VSS2M 52uF
.ends dut
XPcbBuckConverter0 VDD0 VSS0 PcbBuckConverter
Rgnd VSS0 0 0
XPcbModelLumped0 VDD0 VSS0 VDD1 VSS1 PcbModelLumped
Xdut VDD1 VSS1 dut

[['V0', 'VDD0', 'VSS0'], ['V1', 'VDD1', 'VSS1'], ['V1', 'VDD1', 'VSS1'], ['dut.bump.X10Y10X10Y10', 'dut.X10Y10VDD', 'dut.X10Y10VSS'], ['dut.bump.X20Y10X20Y10', 'dut.X20Y10VDD', 'dut.X20Y10VSS'], ['dut.bump.X30Y10X30Y10', 'dut.X30Y10VDD', 'dut.X30Y10VSS'], ['dut.bump.X40Y10X40Y10', 'dut.X40Y10VDD', 'dut.X40Y10VSS'], ['dut.bump.X50Y10X50Y10', 'dut.X50Y10VDD', 'dut.X50Y10VSS'], ['dut.bump.X60Y10X60Y10', 'dut.X60Y10VDD', 'dut.X60Y10VSS'], ['dut.bump.X70Y10X70Y10', 'dut.X70Y10VDD', 'dut.X70Y10VSS'], ['dut.bump.X80Y10X80Y10', 'dut.X80Y10VDD', 'dut.X80Y10VSS'], ['dut.bump.X90Y10X90Y10', 'dut.X90Y10VDD', 'dut.X90Y10VSS'], ['dut.bump.X100Y10X100Y10', 'dut.X100Y10VDD', 'dut.X100Y10VSS'], ['dut.bump.X110Y10X110Y10', 'dut.X110Y10VDD', 'dut.X110Y10VSS'], ['dut.bump.X120Y10X120Y10', 'dut.X120Y10VDD', 'dut.X120Y10VSS'], ['dut.bump.X10Y20X10Y20', 'dut.X10Y20VDD', 'dut.X10Y20VSS'], ['dut.bump.X20Y20X20Y20', 'dut.X20Y20VDD', 'dut.X20Y20VSS'], ['dut.bump.X30Y20X30Y20', 'dut.X30Y20VDD', 'dut.X30Y20VSS'], ['dut.bump.X40Y20X40Y20', 'dut.X40Y20VDD', 'dut.X40Y20VSS'], ['dut.bump.X50Y20X50Y20', 'dut.X50Y20VDD', 'dut.X50Y20VSS'], ['dut.bump.X60Y20X60Y20', 'dut.X60Y20VDD', 'dut.X60Y20VSS'], ['dut.bump.X70Y20X70Y20', 'dut.X70Y20VDD', 'dut.X70Y20VSS'], ['dut.bump.X80Y20X80Y20', 'dut.X80Y20VDD', 'dut.X80Y20VSS'], ['dut.bump.X90Y20X90Y20', 'dut.X90Y20VDD', 'dut.X90Y20VSS'], ['dut.bump.X100Y20X100Y20', 'dut.X100Y20VDD', 'dut.X100Y20VSS'], ['dut.bump.X110Y20X110Y20', 'dut.X110Y20VDD', 'dut.X110Y20VSS'], ['dut.bump.X120Y20X120Y20', 'dut.X120Y20VDD', 'dut.X120Y20VSS'], ['dut.bump.X10Y30X10Y30', 'dut.X10Y30VDD', 'dut.X10Y30VSS'], ['dut.bump.X20Y30X20Y30', 'dut.X20Y30VDD', 'dut.X20Y30VSS'], ['dut.bump.X30Y30X30Y30', 'dut.X30Y30VDD', 'dut.X30Y30VSS'], ['dut.bump.X40Y30X40Y30', 'dut.X40Y30VDD', 'dut.X40Y30VSS'], ['dut.bump.X50Y30X50Y30', 'dut.X50Y30VDD', 'dut.X50Y30VSS'], ['dut.bump.X60Y30X60Y30', 'dut.X60Y30VDD', 'dut.X60Y30VSS'], ['dut.bump.X70Y30X70Y30', 'dut.X70Y30VDD', 'dut.X70Y30VSS'], ['dut.bump.X80Y30X80Y30', 'dut.X80Y30VDD', 'dut.X80Y30VSS'], ['dut.bump.X90Y30X90Y30', 'dut.X90Y30VDD', 'dut.X90Y30VSS'], ['dut.bump.X100Y30X100Y30', 'dut.X100Y30VDD', 'dut.X100Y30VSS'], ['dut.bump.X110Y30X110Y30', 'dut.X110Y30VDD', 'dut.X110Y30VSS'], ['dut.bump.X120Y30X120Y30', 'dut.X120Y30VDD', 'dut.X120Y30VSS'], ['dut.bump.X10Y40X10Y40', 'dut.X10Y40VDD', 'dut.X10Y40VSS'], ['dut.bump.X20Y40X20Y40', 'dut.X20Y40VDD', 'dut.X20Y40VSS'], ['dut.bump.X30Y40X30Y40', 'dut.X30Y40VDD', 'dut.X30Y40VSS'], ['dut.bump.X40Y40X40Y40', 'dut.X40Y40VDD', 'dut.X40Y40VSS'], ['dut.bump.X50Y40X50Y40', 'dut.X50Y40VDD', 'dut.X50Y40VSS'], ['dut.bump.X60Y40X60Y40', 'dut.X60Y40VDD', 'dut.X60Y40VSS'], ['dut.bump.X70Y40X70Y40', 'dut.X70Y40VDD', 'dut.X70Y40VSS'], ['dut.bump.X80Y40X80Y40', 'dut.X80Y40VDD', 'dut.X80Y40VSS'], ['dut.bump.X90Y40X90Y40', 'dut.X90Y40VDD', 'dut.X90Y40VSS'], ['dut.bump.X100Y40X100Y40', 'dut.X100Y40VDD', 'dut.X100Y40VSS'], ['dut.bump.X110Y40X110Y40', 'dut.X110Y40VDD', 'dut.X110Y40VSS'], ['dut.bump.X120Y40X120Y40', 'dut.X120Y40VDD', 'dut.X120Y40VSS'], ['dut.bump.X10Y50X10Y50', 'dut.X10Y50VDD', 'dut.X10Y50VSS'], ['dut.bump.X20Y50X20Y50', 'dut.X20Y50VDD', 'dut.X20Y50VSS'], ['dut.bump.X30Y50X30Y50', 'dut.X30Y50VDD', 'dut.X30Y50VSS'], ['dut.bump.X40Y50X40Y50', 'dut.X40Y50VDD', 'dut.X40Y50VSS'], ['dut.bump.X50Y50X50Y50', 'dut.X50Y50VDD', 'dut.X50Y50VSS'], ['dut.bump.X60Y50X60Y50', 'dut.X60Y50VDD', 'dut.X60Y50VSS'], ['dut.bump.X70Y50X70Y50', 'dut.X70Y50VDD', 'dut.X70Y50VSS'], ['dut.bump.X80Y50X80Y50', 'dut.X80Y50VDD', 'dut.X80Y50VSS'], ['dut.bump.X90Y50X90Y50', 'dut.X90Y50VDD', 'dut.X90Y50VSS'], ['dut.bump.X100Y50X100Y50', 'dut.X100Y50VDD', 'dut.X100Y50VSS'], ['dut.bump.X110Y50X110Y50', 'dut.X110Y50VDD', 'dut.X110Y50VSS'], ['dut.bump.X120Y50X120Y50', 'dut.X120Y50VDD', 'dut.X120Y50VSS'], ['dut.bump.X10Y60X10Y60', 'dut.X10Y60VDD', 'dut.X10Y60VSS'], ['dut.bump.X20Y60X20Y60', 'dut.X20Y60VDD', 'dut.X20Y60VSS'], ['dut.bump.X30Y60X30Y60', 'dut.X30Y60VDD', 'dut.X30Y60VSS'], ['dut.bump.X40Y60X40Y60', 'dut.X40Y60VDD', 'dut.X40Y60VSS'], ['dut.bump.X50Y60X50Y60', 'dut.X50Y60VDD', 'dut.X50Y60VSS'], ['dut.bump.X60Y60X60Y60', 'dut.X60Y60VDD', 'dut.X60Y60VSS'], ['dut.bump.X70Y60X70Y60', 'dut.X70Y60VDD', 'dut.X70Y60VSS'], ['dut.bump.X80Y60X80Y60', 'dut.X80Y60VDD', 'dut.X80Y60VSS'], ['dut.bump.X90Y60X90Y60', 'dut.X90Y60VDD', 'dut.X90Y60VSS'], ['dut.bump.X100Y60X100Y60', 'dut.X100Y60VDD', 'dut.X100Y60VSS'], ['dut.bump.X110Y60X110Y60', 'dut.X110Y60VDD', 'dut.X110Y60VSS'], ['dut.bump.X120Y60X120Y60', 'dut.X120Y60VDD', 'dut.X120Y60VSS'], ['dut.bump.X10Y70X10Y70', 'dut.X10Y70VDD', 'dut.X10Y70VSS'], ['dut.bump.X20Y70X20Y70', 'dut.X20Y70VDD', 'dut.X20Y70VSS'], ['dut.bump.X30Y70X30Y70', 'dut.X30Y70VDD', 'dut.X30Y70VSS'], ['dut.bump.X40Y70X40Y70', 'dut.X40Y70VDD', 'dut.X40Y70VSS'], ['dut.bump.X50Y70X50Y70', 'dut.X50Y70VDD', 'dut.X50Y70VSS'], ['dut.bump.X60Y70X60Y70', 'dut.X60Y70VDD', 'dut.X60Y70VSS'], ['dut.bump.X70Y70X70Y70', 'dut.X70Y70VDD', 'dut.X70Y70VSS'], ['dut.bump.X80Y70X80Y70', 'dut.X80Y70VDD', 'dut.X80Y70VSS'], ['dut.bump.X90Y70X90Y70', 'dut.X90Y70VDD', 'dut.X90Y70VSS'], ['dut.bump.X100Y70X100Y70', 'dut.X100Y70VDD', 'dut.X100Y70VSS'], ['dut.bump.X110Y70X110Y70', 'dut.X110Y70VDD', 'dut.X110Y70VSS'], ['dut.bump.X120Y70X120Y70', 'dut.X120Y70VDD', 'dut.X120Y70VSS'], ['dut.bump.X10Y80X10Y80', 'dut.X10Y80VDD', 'dut.X10Y80VSS'], ['dut.bump.X20Y80X20Y80', 'dut.X20Y80VDD', 'dut.X20Y80VSS'], ['dut.bump.X30Y80X30Y80', 'dut.X30Y80VDD', 'dut.X30Y80VSS'], ['dut.bump.X40Y80X40Y80', 'dut.X40Y80VDD', 'dut.X40Y80VSS'], ['dut.bump.X50Y80X50Y80', 'dut.X50Y80VDD', 'dut.X50Y80VSS'], ['dut.bump.X60Y80X60Y80', 'dut.X60Y80VDD', 'dut.X60Y80VSS'], ['dut.bump.X70Y80X70Y80', 'dut.X70Y80VDD', 'dut.X70Y80VSS'], ['dut.bump.X80Y80X80Y80', 'dut.X80Y80VDD', 'dut.X80Y80VSS'], ['dut.bump.X90Y80X90Y80', 'dut.X90Y80VDD', 'dut.X90Y80VSS'], ['dut.bump.X100Y80X100Y80', 'dut.X100Y80VDD', 'dut.X100Y80VSS'], ['dut.bump.X110Y80X110Y80', 'dut.X110Y80VDD', 'dut.X110Y80VSS'], ['dut.bump.X120Y80X120Y80', 'dut.X120Y80VDD', 'dut.X120Y80VSS'], ['dut.bump.X10Y90X10Y90', 'dut.X10Y90VDD', 'dut.X10Y90VSS'], ['dut.bump.X20Y90X20Y90', 'dut.X20Y90VDD', 'dut.X20Y90VSS'], ['dut.bump.X30Y90X30Y90', 'dut.X30Y90VDD', 'dut.X30Y90VSS'], ['dut.bump.X40Y90X40Y90', 'dut.X40Y90VDD', 'dut.X40Y90VSS'], ['dut.bump.X50Y90X50Y90', 'dut.X50Y90VDD', 'dut.X50Y90VSS'], ['dut.bump.X60Y90X60Y90', 'dut.X60Y90VDD', 'dut.X60Y90VSS'], ['dut.bump.X70Y90X70Y90', 'dut.X70Y90VDD', 'dut.X70Y90VSS'], ['dut.bump.X80Y90X80Y90', 'dut.X80Y90VDD', 'dut.X80Y90VSS'], ['dut.bump.X90Y90X90Y90', 'dut.X90Y90VDD', 'dut.X90Y90VSS'], ['dut.bump.X100Y90X100Y90', 'dut.X100Y90VDD', 'dut.X100Y90VSS'], ['dut.bump.X110Y90X110Y90', 'dut.X110Y90VDD', 'dut.X110Y90VSS'], ['dut.bump.X120Y90X120Y90', 'dut.X120Y90VDD', 'dut.X120Y90VSS'], ['dut.bump.X10Y100X10Y100', 'dut.X10Y100VDD', 'dut.X10Y100VSS'], ['dut.bump.X20Y100X20Y100', 'dut.X20Y100VDD', 'dut.X20Y100VSS'], ['dut.bump.X30Y100X30Y100', 'dut.X30Y100VDD', 'dut.X30Y100VSS'], ['dut.bump.X40Y100X40Y100', 'dut.X40Y100VDD', 'dut.X40Y100VSS'], ['dut.bump.X50Y100X50Y100', 'dut.X50Y100VDD', 'dut.X50Y100VSS'], ['dut.bump.X60Y100X60Y100', 'dut.X60Y100VDD', 'dut.X60Y100VSS'], ['dut.bump.X70Y100X70Y100', 'dut.X70Y100VDD', 'dut.X70Y100VSS'], ['dut.bump.X80Y100X80Y100', 'dut.X80Y100VDD', 'dut.X80Y100VSS'], ['dut.bump.X90Y100X90Y100', 'dut.X90Y100VDD', 'dut.X90Y100VSS'], ['dut.bump.X100Y100X100Y100', 'dut.X100Y100VDD', 'dut.X100Y100VSS'], ['dut.bump.X110Y100X110Y100', 'dut.X110Y100VDD', 'dut.X110Y100VSS'], ['dut.bump.X120Y100X120Y100', 'dut.X120Y100VDD', 'dut.X120Y100VSS'], ['dut.bump.X10Y110X10Y110', 'dut.X10Y110VDD', 'dut.X10Y110VSS'], ['dut.bump.X20Y110X20Y110', 'dut.X20Y110VDD', 'dut.X20Y110VSS'], ['dut.bump.X30Y110X30Y110', 'dut.X30Y110VDD', 'dut.X30Y110VSS'], ['dut.bump.X40Y110X40Y110', 'dut.X40Y110VDD', 'dut.X40Y110VSS'], ['dut.bump.X50Y110X50Y110', 'dut.X50Y110VDD', 'dut.X50Y110VSS'], ['dut.bump.X60Y110X60Y110', 'dut.X60Y110VDD', 'dut.X60Y110VSS'], ['dut.bump.X70Y110X70Y110', 'dut.X70Y110VDD', 'dut.X70Y110VSS'], ['dut.bump.X80Y110X80Y110', 'dut.X80Y110VDD', 'dut.X80Y110VSS'], ['dut.bump.X90Y110X90Y110', 'dut.X90Y110VDD', 'dut.X90Y110VSS'], ['dut.bump.X100Y110X100Y110', 'dut.X100Y110VDD', 'dut.X100Y110VSS'], ['dut.bump.X110Y110X110Y110', 'dut.X110Y110VDD', 'dut.X110Y110VSS'], ['dut.bump.X120Y110X120Y110', 'dut.X120Y110VDD', 'dut.X120Y110VSS'], ['dut.bump.X10Y120X10Y120', 'dut.X10Y120VDD', 'dut.X10Y120VSS'], ['dut.bump.X20Y120X20Y120', 'dut.X20Y120VDD', 'dut.X20Y120VSS'], ['dut.bump.X30Y120X30Y120', 'dut.X30Y120VDD', 'dut.X30Y120VSS'], ['dut.bump.X40Y120X40Y120', 'dut.X40Y120VDD', 'dut.X40Y120VSS'], ['dut.bump.X50Y120X50Y120', 'dut.X50Y120VDD', 'dut.X50Y120VSS'], ['dut.bump.X60Y120X60Y120', 'dut.X60Y120VDD', 'dut.X60Y120VSS'], ['dut.bump.X70Y120X70Y120', 'dut.X70Y120VDD', 'dut.X70Y120VSS'], ['dut.bump.X80Y120X80Y120', 'dut.X80Y120VDD', 'dut.X80Y120VSS'], ['dut.bump.X90Y120X90Y120', 'dut.X90Y120VDD', 'dut.X90Y120VSS'], ['dut.bump.X100Y120X100Y120', 'dut.X100Y120VDD', 'dut.X100Y120VSS'], ['dut.bump.X110Y120X110Y120', 'dut.X110Y120VDD', 'dut.X110Y120VSS'], ['dut.bump.X120Y120X120Y120', 'dut.X120Y120VDD', 'dut.X120Y120VSS']]
.title 20200622-105341
.option rshunt = 1.0e12
.subckt Regulator VDD VSS
Vs VDD VSS 1.1
.ends Regulator

.subckt ChipPackage VDD1 VSS1 VDD2 VSS2
RsVDD VDD1 VDDMS 0.55mOhm
LsVDD VDDMS VDD2 0.06nH
RsVSS VSS1 VSSMS 0.55mOhm
LsVSS VSSMS VSS2 0.06nH
Rp VDD2 VDD2M 0.1mOhm
Lp VSS2 VSS2M 0.0028nH
Cp VDD2M VSS2M 52uF
.ends ChipPackage

.subckt ChipBump VDD1 VSS1 VDD2 VSS2
RX0Y0VDD VDD1 X0Y0VDDM 20mOhm
LX0Y0VDD X0Y0VDDM VDD2 0.036nH
RX0Y0VSS VSS1 X0Y0VSSM 20mOhm
LX0Y0VSS X0Y0VSSM VSS2 0.036nH
RX0Y1VDD VDD1 X0Y1VDDM 20mOhm
LX0Y1VDD X0Y1VDDM VDD2 0.036nH
RX0Y1VSS VSS1 X0Y1VSSM 20mOhm
LX0Y1VSS X0Y1VSSM VSS2 0.036nH
RX0Y2VDD VDD1 X0Y2VDDM 20mOhm
LX0Y2VDD X0Y2VDDM VDD2 0.036nH
RX0Y2VSS VSS1 X0Y2VSSM 20mOhm
LX0Y2VSS X0Y2VSSM VSS2 0.036nH
RX0Y3VDD VDD1 X0Y3VDDM 20mOhm
LX0Y3VDD X0Y3VDDM VDD2 0.036nH
RX0Y3VSS VSS1 X0Y3VSSM 20mOhm
LX0Y3VSS X0Y3VSSM VSS2 0.036nH
RX0Y4VDD VDD1 X0Y4VDDM 20mOhm
LX0Y4VDD X0Y4VDDM VDD2 0.036nH
RX0Y4VSS VSS1 X0Y4VSSM 20mOhm
LX0Y4VSS X0Y4VSSM VSS2 0.036nH
RX0Y5VDD VDD1 X0Y5VDDM 20mOhm
LX0Y5VDD X0Y5VDDM VDD2 0.036nH
RX0Y5VSS VSS1 X0Y5VSSM 20mOhm
LX0Y5VSS X0Y5VSSM VSS2 0.036nH
RX0Y6VDD VDD1 X0Y6VDDM 20mOhm
LX0Y6VDD X0Y6VDDM VDD2 0.036nH
RX0Y6VSS VSS1 X0Y6VSSM 20mOhm
LX0Y6VSS X0Y6VSSM VSS2 0.036nH
RX0Y7VDD VDD1 X0Y7VDDM 20mOhm
LX0Y7VDD X0Y7VDDM VDD2 0.036nH
RX0Y7VSS VSS1 X0Y7VSSM 20mOhm
LX0Y7VSS X0Y7VSSM VSS2 0.036nH
RX0Y8VDD VDD1 X0Y8VDDM 20mOhm
LX0Y8VDD X0Y8VDDM VDD2 0.036nH
RX0Y8VSS VSS1 X0Y8VSSM 20mOhm
LX0Y8VSS X0Y8VSSM VSS2 0.036nH
RX0Y9VDD VDD1 X0Y9VDDM 20mOhm
LX0Y9VDD X0Y9VDDM VDD2 0.036nH
RX0Y9VSS VSS1 X0Y9VSSM 20mOhm
LX0Y9VSS X0Y9VSSM VSS2 0.036nH
RX0Y10VDD VDD1 X0Y10VDDM 20mOhm
LX0Y10VDD X0Y10VDDM VDD2 0.036nH
RX0Y10VSS VSS1 X0Y10VSSM 20mOhm
LX0Y10VSS X0Y10VSSM VSS2 0.036nH
RX0Y11VDD VDD1 X0Y11VDDM 20mOhm
LX0Y11VDD X0Y11VDDM VDD2 0.036nH
RX0Y11VSS VSS1 X0Y11VSSM 20mOhm
LX0Y11VSS X0Y11VSSM VSS2 0.036nH
RX1Y0VDD VDD1 X1Y0VDDM 20mOhm
LX1Y0VDD X1Y0VDDM VDD2 0.036nH
RX1Y0VSS VSS1 X1Y0VSSM 20mOhm
LX1Y0VSS X1Y0VSSM VSS2 0.036nH
RX1Y1VDD VDD1 X1Y1VDDM 20mOhm
LX1Y1VDD X1Y1VDDM VDD2 0.036nH
RX1Y1VSS VSS1 X1Y1VSSM 20mOhm
LX1Y1VSS X1Y1VSSM VSS2 0.036nH
RX1Y2VDD VDD1 X1Y2VDDM 20mOhm
LX1Y2VDD X1Y2VDDM VDD2 0.036nH
RX1Y2VSS VSS1 X1Y2VSSM 20mOhm
LX1Y2VSS X1Y2VSSM VSS2 0.036nH
RX1Y3VDD VDD1 X1Y3VDDM 20mOhm
LX1Y3VDD X1Y3VDDM VDD2 0.036nH
RX1Y3VSS VSS1 X1Y3VSSM 20mOhm
LX1Y3VSS X1Y3VSSM VSS2 0.036nH
RX1Y4VDD VDD1 X1Y4VDDM 20mOhm
LX1Y4VDD X1Y4VDDM VDD2 0.036nH
RX1Y4VSS VSS1 X1Y4VSSM 20mOhm
LX1Y4VSS X1Y4VSSM VSS2 0.036nH
RX1Y5VDD VDD1 X1Y5VDDM 20mOhm
LX1Y5VDD X1Y5VDDM VDD2 0.036nH
RX1Y5VSS VSS1 X1Y5VSSM 20mOhm
LX1Y5VSS X1Y5VSSM VSS2 0.036nH
RX1Y6VDD VDD1 X1Y6VDDM 20mOhm
LX1Y6VDD X1Y6VDDM VDD2 0.036nH
RX1Y6VSS VSS1 X1Y6VSSM 20mOhm
LX1Y6VSS X1Y6VSSM VSS2 0.036nH
RX1Y7VDD VDD1 X1Y7VDDM 20mOhm
LX1Y7VDD X1Y7VDDM VDD2 0.036nH
RX1Y7VSS VSS1 X1Y7VSSM 20mOhm
LX1Y7VSS X1Y7VSSM VSS2 0.036nH
RX1Y8VDD VDD1 X1Y8VDDM 20mOhm
LX1Y8VDD X1Y8VDDM VDD2 0.036nH
RX1Y8VSS VSS1 X1Y8VSSM 20mOhm
LX1Y8VSS X1Y8VSSM VSS2 0.036nH
RX1Y9VDD VDD1 X1Y9VDDM 20mOhm
LX1Y9VDD X1Y9VDDM VDD2 0.036nH
RX1Y9VSS VSS1 X1Y9VSSM 20mOhm
LX1Y9VSS X1Y9VSSM VSS2 0.036nH
RX1Y10VDD VDD1 X1Y10VDDM 20mOhm
LX1Y10VDD X1Y10VDDM VDD2 0.036nH
RX1Y10VSS VSS1 X1Y10VSSM 20mOhm
LX1Y10VSS X1Y10VSSM VSS2 0.036nH
RX1Y11VDD VDD1 X1Y11VDDM 20mOhm
LX1Y11VDD X1Y11VDDM VDD2 0.036nH
RX1Y11VSS VSS1 X1Y11VSSM 20mOhm
LX1Y11VSS X1Y11VSSM VSS2 0.036nH
RX2Y0VDD VDD1 X2Y0VDDM 20mOhm
LX2Y0VDD X2Y0VDDM VDD2 0.036nH
RX2Y0VSS VSS1 X2Y0VSSM 20mOhm
LX2Y0VSS X2Y0VSSM VSS2 0.036nH
RX2Y1VDD VDD1 X2Y1VDDM 20mOhm
LX2Y1VDD X2Y1VDDM VDD2 0.036nH
RX2Y1VSS VSS1 X2Y1VSSM 20mOhm
LX2Y1VSS X2Y1VSSM VSS2 0.036nH
RX2Y2VDD VDD1 X2Y2VDDM 20mOhm
LX2Y2VDD X2Y2VDDM VDD2 0.036nH
RX2Y2VSS VSS1 X2Y2VSSM 20mOhm
LX2Y2VSS X2Y2VSSM VSS2 0.036nH
RX2Y3VDD VDD1 X2Y3VDDM 20mOhm
LX2Y3VDD X2Y3VDDM VDD2 0.036nH
RX2Y3VSS VSS1 X2Y3VSSM 20mOhm
LX2Y3VSS X2Y3VSSM VSS2 0.036nH
RX2Y4VDD VDD1 X2Y4VDDM 20mOhm
LX2Y4VDD X2Y4VDDM VDD2 0.036nH
RX2Y4VSS VSS1 X2Y4VSSM 20mOhm
LX2Y4VSS X2Y4VSSM VSS2 0.036nH
RX2Y5VDD VDD1 X2Y5VDDM 20mOhm
LX2Y5VDD X2Y5VDDM VDD2 0.036nH
RX2Y5VSS VSS1 X2Y5VSSM 20mOhm
LX2Y5VSS X2Y5VSSM VSS2 0.036nH
RX2Y6VDD VDD1 X2Y6VDDM 20mOhm
LX2Y6VDD X2Y6VDDM VDD2 0.036nH
RX2Y6VSS VSS1 X2Y6VSSM 20mOhm
LX2Y6VSS X2Y6VSSM VSS2 0.036nH
RX2Y7VDD VDD1 X2Y7VDDM 20mOhm
LX2Y7VDD X2Y7VDDM VDD2 0.036nH
RX2Y7VSS VSS1 X2Y7VSSM 20mOhm
LX2Y7VSS X2Y7VSSM VSS2 0.036nH
RX2Y8VDD VDD1 X2Y8VDDM 20mOhm
LX2Y8VDD X2Y8VDDM VDD2 0.036nH
RX2Y8VSS VSS1 X2Y8VSSM 20mOhm
LX2Y8VSS X2Y8VSSM VSS2 0.036nH
RX2Y9VDD VDD1 X2Y9VDDM 20mOhm
LX2Y9VDD X2Y9VDDM VDD2 0.036nH
RX2Y9VSS VSS1 X2Y9VSSM 20mOhm
LX2Y9VSS X2Y9VSSM VSS2 0.036nH
RX2Y10VDD VDD1 X2Y10VDDM 20mOhm
LX2Y10VDD X2Y10VDDM VDD2 0.036nH
RX2Y10VSS VSS1 X2Y10VSSM 20mOhm
LX2Y10VSS X2Y10VSSM VSS2 0.036nH
RX2Y11VDD VDD1 X2Y11VDDM 20mOhm
LX2Y11VDD X2Y11VDDM VDD2 0.036nH
RX2Y11VSS VSS1 X2Y11VSSM 20mOhm
LX2Y11VSS X2Y11VSSM VSS2 0.036nH
RX3Y0VDD VDD1 X3Y0VDDM 20mOhm
LX3Y0VDD X3Y0VDDM VDD2 0.036nH
RX3Y0VSS VSS1 X3Y0VSSM 20mOhm
LX3Y0VSS X3Y0VSSM VSS2 0.036nH
RX3Y1VDD VDD1 X3Y1VDDM 20mOhm
LX3Y1VDD X3Y1VDDM VDD2 0.036nH
RX3Y1VSS VSS1 X3Y1VSSM 20mOhm
LX3Y1VSS X3Y1VSSM VSS2 0.036nH
RX3Y2VDD VDD1 X3Y2VDDM 20mOhm
LX3Y2VDD X3Y2VDDM VDD2 0.036nH
RX3Y2VSS VSS1 X3Y2VSSM 20mOhm
LX3Y2VSS X3Y2VSSM VSS2 0.036nH
RX3Y3VDD VDD1 X3Y3VDDM 20mOhm
LX3Y3VDD X3Y3VDDM VDD2 0.036nH
RX3Y3VSS VSS1 X3Y3VSSM 20mOhm
LX3Y3VSS X3Y3VSSM VSS2 0.036nH
RX3Y4VDD VDD1 X3Y4VDDM 20mOhm
LX3Y4VDD X3Y4VDDM VDD2 0.036nH
RX3Y4VSS VSS1 X3Y4VSSM 20mOhm
LX3Y4VSS X3Y4VSSM VSS2 0.036nH
RX3Y5VDD VDD1 X3Y5VDDM 20mOhm
LX3Y5VDD X3Y5VDDM VDD2 0.036nH
RX3Y5VSS VSS1 X3Y5VSSM 20mOhm
LX3Y5VSS X3Y5VSSM VSS2 0.036nH
RX3Y6VDD VDD1 X3Y6VDDM 20mOhm
LX3Y6VDD X3Y6VDDM VDD2 0.036nH
RX3Y6VSS VSS1 X3Y6VSSM 20mOhm
LX3Y6VSS X3Y6VSSM VSS2 0.036nH
RX3Y7VDD VDD1 X3Y7VDDM 20mOhm
LX3Y7VDD X3Y7VDDM VDD2 0.036nH
RX3Y7VSS VSS1 X3Y7VSSM 20mOhm
LX3Y7VSS X3Y7VSSM VSS2 0.036nH
RX3Y8VDD VDD1 X3Y8VDDM 20mOhm
LX3Y8VDD X3Y8VDDM VDD2 0.036nH
RX3Y8VSS VSS1 X3Y8VSSM 20mOhm
LX3Y8VSS X3Y8VSSM VSS2 0.036nH
RX3Y9VDD VDD1 X3Y9VDDM 20mOhm
LX3Y9VDD X3Y9VDDM VDD2 0.036nH
RX3Y9VSS VSS1 X3Y9VSSM 20mOhm
LX3Y9VSS X3Y9VSSM VSS2 0.036nH
RX3Y10VDD VDD1 X3Y10VDDM 20mOhm
LX3Y10VDD X3Y10VDDM VDD2 0.036nH
RX3Y10VSS VSS1 X3Y10VSSM 20mOhm
LX3Y10VSS X3Y10VSSM VSS2 0.036nH
RX3Y11VDD VDD1 X3Y11VDDM 20mOhm
LX3Y11VDD X3Y11VDDM VDD2 0.036nH
RX3Y11VSS VSS1 X3Y11VSSM 20mOhm
LX3Y11VSS X3Y11VSSM VSS2 0.036nH
RX4Y0VDD VDD1 X4Y0VDDM 20mOhm
LX4Y0VDD X4Y0VDDM VDD2 0.036nH
RX4Y0VSS VSS1 X4Y0VSSM 20mOhm
LX4Y0VSS X4Y0VSSM VSS2 0.036nH
RX4Y1VDD VDD1 X4Y1VDDM 20mOhm
LX4Y1VDD X4Y1VDDM VDD2 0.036nH
RX4Y1VSS VSS1 X4Y1VSSM 20mOhm
LX4Y1VSS X4Y1VSSM VSS2 0.036nH
RX4Y2VDD VDD1 X4Y2VDDM 20mOhm
LX4Y2VDD X4Y2VDDM VDD2 0.036nH
RX4Y2VSS VSS1 X4Y2VSSM 20mOhm
LX4Y2VSS X4Y2VSSM VSS2 0.036nH
RX4Y3VDD VDD1 X4Y3VDDM 20mOhm
LX4Y3VDD X4Y3VDDM VDD2 0.036nH
RX4Y3VSS VSS1 X4Y3VSSM 20mOhm
LX4Y3VSS X4Y3VSSM VSS2 0.036nH
RX4Y4VDD VDD1 X4Y4VDDM 20mOhm
LX4Y4VDD X4Y4VDDM VDD2 0.036nH
RX4Y4VSS VSS1 X4Y4VSSM 20mOhm
LX4Y4VSS X4Y4VSSM VSS2 0.036nH
RX4Y5VDD VDD1 X4Y5VDDM 20mOhm
LX4Y5VDD X4Y5VDDM VDD2 0.036nH
RX4Y5VSS VSS1 X4Y5VSSM 20mOhm
LX4Y5VSS X4Y5VSSM VSS2 0.036nH
RX4Y6VDD VDD1 X4Y6VDDM 20mOhm
LX4Y6VDD X4Y6VDDM VDD2 0.036nH
RX4Y6VSS VSS1 X4Y6VSSM 20mOhm
LX4Y6VSS X4Y6VSSM VSS2 0.036nH
RX4Y7VDD VDD1 X4Y7VDDM 20mOhm
LX4Y7VDD X4Y7VDDM VDD2 0.036nH
RX4Y7VSS VSS1 X4Y7VSSM 20mOhm
LX4Y7VSS X4Y7VSSM VSS2 0.036nH
RX4Y8VDD VDD1 X4Y8VDDM 20mOhm
LX4Y8VDD X4Y8VDDM VDD2 0.036nH
RX4Y8VSS VSS1 X4Y8VSSM 20mOhm
LX4Y8VSS X4Y8VSSM VSS2 0.036nH
RX4Y9VDD VDD1 X4Y9VDDM 20mOhm
LX4Y9VDD X4Y9VDDM VDD2 0.036nH
RX4Y9VSS VSS1 X4Y9VSSM 20mOhm
LX4Y9VSS X4Y9VSSM VSS2 0.036nH
RX4Y10VDD VDD1 X4Y10VDDM 20mOhm
LX4Y10VDD X4Y10VDDM VDD2 0.036nH
RX4Y10VSS VSS1 X4Y10VSSM 20mOhm
LX4Y10VSS X4Y10VSSM VSS2 0.036nH
RX4Y11VDD VDD1 X4Y11VDDM 20mOhm
LX4Y11VDD X4Y11VDDM VDD2 0.036nH
RX4Y11VSS VSS1 X4Y11VSSM 20mOhm
LX4Y11VSS X4Y11VSSM VSS2 0.036nH
RX5Y0VDD VDD1 X5Y0VDDM 20mOhm
LX5Y0VDD X5Y0VDDM VDD2 0.036nH
RX5Y0VSS VSS1 X5Y0VSSM 20mOhm
LX5Y0VSS X5Y0VSSM VSS2 0.036nH
RX5Y1VDD VDD1 X5Y1VDDM 20mOhm
LX5Y1VDD X5Y1VDDM VDD2 0.036nH
RX5Y1VSS VSS1 X5Y1VSSM 20mOhm
LX5Y1VSS X5Y1VSSM VSS2 0.036nH
RX5Y2VDD VDD1 X5Y2VDDM 20mOhm
LX5Y2VDD X5Y2VDDM VDD2 0.036nH
RX5Y2VSS VSS1 X5Y2VSSM 20mOhm
LX5Y2VSS X5Y2VSSM VSS2 0.036nH
RX5Y3VDD VDD1 X5Y3VDDM 20mOhm
LX5Y3VDD X5Y3VDDM VDD2 0.036nH
RX5Y3VSS VSS1 X5Y3VSSM 20mOhm
LX5Y3VSS X5Y3VSSM VSS2 0.036nH
RX5Y4VDD VDD1 X5Y4VDDM 20mOhm
LX5Y4VDD X5Y4VDDM VDD2 0.036nH
RX5Y4VSS VSS1 X5Y4VSSM 20mOhm
LX5Y4VSS X5Y4VSSM VSS2 0.036nH
RX5Y5VDD VDD1 X5Y5VDDM 20mOhm
LX5Y5VDD X5Y5VDDM VDD2 0.036nH
RX5Y5VSS VSS1 X5Y5VSSM 20mOhm
LX5Y5VSS X5Y5VSSM VSS2 0.036nH
RX5Y6VDD VDD1 X5Y6VDDM 20mOhm
LX5Y6VDD X5Y6VDDM VDD2 0.036nH
RX5Y6VSS VSS1 X5Y6VSSM 20mOhm
LX5Y6VSS X5Y6VSSM VSS2 0.036nH
RX5Y7VDD VDD1 X5Y7VDDM 20mOhm
LX5Y7VDD X5Y7VDDM VDD2 0.036nH
RX5Y7VSS VSS1 X5Y7VSSM 20mOhm
LX5Y7VSS X5Y7VSSM VSS2 0.036nH
RX5Y8VDD VDD1 X5Y8VDDM 20mOhm
LX5Y8VDD X5Y8VDDM VDD2 0.036nH
RX5Y8VSS VSS1 X5Y8VSSM 20mOhm
LX5Y8VSS X5Y8VSSM VSS2 0.036nH
RX5Y9VDD VDD1 X5Y9VDDM 20mOhm
LX5Y9VDD X5Y9VDDM VDD2 0.036nH
RX5Y9VSS VSS1 X5Y9VSSM 20mOhm
LX5Y9VSS X5Y9VSSM VSS2 0.036nH
RX5Y10VDD VDD1 X5Y10VDDM 20mOhm
LX5Y10VDD X5Y10VDDM VDD2 0.036nH
RX5Y10VSS VSS1 X5Y10VSSM 20mOhm
LX5Y10VSS X5Y10VSSM VSS2 0.036nH
RX5Y11VDD VDD1 X5Y11VDDM 20mOhm
LX5Y11VDD X5Y11VDDM VDD2 0.036nH
RX5Y11VSS VSS1 X5Y11VSSM 20mOhm
LX5Y11VSS X5Y11VSSM VSS2 0.036nH
RX6Y0VDD VDD1 X6Y0VDDM 20mOhm
LX6Y0VDD X6Y0VDDM VDD2 0.036nH
RX6Y0VSS VSS1 X6Y0VSSM 20mOhm
LX6Y0VSS X6Y0VSSM VSS2 0.036nH
RX6Y1VDD VDD1 X6Y1VDDM 20mOhm
LX6Y1VDD X6Y1VDDM VDD2 0.036nH
RX6Y1VSS VSS1 X6Y1VSSM 20mOhm
LX6Y1VSS X6Y1VSSM VSS2 0.036nH
RX6Y2VDD VDD1 X6Y2VDDM 20mOhm
LX6Y2VDD X6Y2VDDM VDD2 0.036nH
RX6Y2VSS VSS1 X6Y2VSSM 20mOhm
LX6Y2VSS X6Y2VSSM VSS2 0.036nH
RX6Y3VDD VDD1 X6Y3VDDM 20mOhm
LX6Y3VDD X6Y3VDDM VDD2 0.036nH
RX6Y3VSS VSS1 X6Y3VSSM 20mOhm
LX6Y3VSS X6Y3VSSM VSS2 0.036nH
RX6Y4VDD VDD1 X6Y4VDDM 20mOhm
LX6Y4VDD X6Y4VDDM VDD2 0.036nH
RX6Y4VSS VSS1 X6Y4VSSM 20mOhm
LX6Y4VSS X6Y4VSSM VSS2 0.036nH
RX6Y5VDD VDD1 X6Y5VDDM 20mOhm
LX6Y5VDD X6Y5VDDM VDD2 0.036nH
RX6Y5VSS VSS1 X6Y5VSSM 20mOhm
LX6Y5VSS X6Y5VSSM VSS2 0.036nH
RX6Y6VDD VDD1 X6Y6VDDM 20mOhm
LX6Y6VDD X6Y6VDDM VDD2 0.036nH
RX6Y6VSS VSS1 X6Y6VSSM 20mOhm
LX6Y6VSS X6Y6VSSM VSS2 0.036nH
RX6Y7VDD VDD1 X6Y7VDDM 20mOhm
LX6Y7VDD X6Y7VDDM VDD2 0.036nH
RX6Y7VSS VSS1 X6Y7VSSM 20mOhm
LX6Y7VSS X6Y7VSSM VSS2 0.036nH
RX6Y8VDD VDD1 X6Y8VDDM 20mOhm
LX6Y8VDD X6Y8VDDM VDD2 0.036nH
RX6Y8VSS VSS1 X6Y8VSSM 20mOhm
LX6Y8VSS X6Y8VSSM VSS2 0.036nH
RX6Y9VDD VDD1 X6Y9VDDM 20mOhm
LX6Y9VDD X6Y9VDDM VDD2 0.036nH
RX6Y9VSS VSS1 X6Y9VSSM 20mOhm
LX6Y9VSS X6Y9VSSM VSS2 0.036nH
RX6Y10VDD VDD1 X6Y10VDDM 20mOhm
LX6Y10VDD X6Y10VDDM VDD2 0.036nH
RX6Y10VSS VSS1 X6Y10VSSM 20mOhm
LX6Y10VSS X6Y10VSSM VSS2 0.036nH
RX6Y11VDD VDD1 X6Y11VDDM 20mOhm
LX6Y11VDD X6Y11VDDM VDD2 0.036nH
RX6Y11VSS VSS1 X6Y11VSSM 20mOhm
LX6Y11VSS X6Y11VSSM VSS2 0.036nH
RX7Y0VDD VDD1 X7Y0VDDM 20mOhm
LX7Y0VDD X7Y0VDDM VDD2 0.036nH
RX7Y0VSS VSS1 X7Y0VSSM 20mOhm
LX7Y0VSS X7Y0VSSM VSS2 0.036nH
RX7Y1VDD VDD1 X7Y1VDDM 20mOhm
LX7Y1VDD X7Y1VDDM VDD2 0.036nH
RX7Y1VSS VSS1 X7Y1VSSM 20mOhm
LX7Y1VSS X7Y1VSSM VSS2 0.036nH
RX7Y2VDD VDD1 X7Y2VDDM 20mOhm
LX7Y2VDD X7Y2VDDM VDD2 0.036nH
RX7Y2VSS VSS1 X7Y2VSSM 20mOhm
LX7Y2VSS X7Y2VSSM VSS2 0.036nH
RX7Y3VDD VDD1 X7Y3VDDM 20mOhm
LX7Y3VDD X7Y3VDDM VDD2 0.036nH
RX7Y3VSS VSS1 X7Y3VSSM 20mOhm
LX7Y3VSS X7Y3VSSM VSS2 0.036nH
RX7Y4VDD VDD1 X7Y4VDDM 20mOhm
LX7Y4VDD X7Y4VDDM VDD2 0.036nH
RX7Y4VSS VSS1 X7Y4VSSM 20mOhm
LX7Y4VSS X7Y4VSSM VSS2 0.036nH
RX7Y5VDD VDD1 X7Y5VDDM 20mOhm
LX7Y5VDD X7Y5VDDM VDD2 0.036nH
RX7Y5VSS VSS1 X7Y5VSSM 20mOhm
LX7Y5VSS X7Y5VSSM VSS2 0.036nH
RX7Y6VDD VDD1 X7Y6VDDM 20mOhm
LX7Y6VDD X7Y6VDDM VDD2 0.036nH
RX7Y6VSS VSS1 X7Y6VSSM 20mOhm
LX7Y6VSS X7Y6VSSM VSS2 0.036nH
RX7Y7VDD VDD1 X7Y7VDDM 20mOhm
LX7Y7VDD X7Y7VDDM VDD2 0.036nH
RX7Y7VSS VSS1 X7Y7VSSM 20mOhm
LX7Y7VSS X7Y7VSSM VSS2 0.036nH
RX7Y8VDD VDD1 X7Y8VDDM 20mOhm
LX7Y8VDD X7Y8VDDM VDD2 0.036nH
RX7Y8VSS VSS1 X7Y8VSSM 20mOhm
LX7Y8VSS X7Y8VSSM VSS2 0.036nH
RX7Y9VDD VDD1 X7Y9VDDM 20mOhm
LX7Y9VDD X7Y9VDDM VDD2 0.036nH
RX7Y9VSS VSS1 X7Y9VSSM 20mOhm
LX7Y9VSS X7Y9VSSM VSS2 0.036nH
RX7Y10VDD VDD1 X7Y10VDDM 20mOhm
LX7Y10VDD X7Y10VDDM VDD2 0.036nH
RX7Y10VSS VSS1 X7Y10VSSM 20mOhm
LX7Y10VSS X7Y10VSSM VSS2 0.036nH
RX7Y11VDD VDD1 X7Y11VDDM 20mOhm
LX7Y11VDD X7Y11VDDM VDD2 0.036nH
RX7Y11VSS VSS1 X7Y11VSSM 20mOhm
LX7Y11VSS X7Y11VSSM VSS2 0.036nH
RX8Y0VDD VDD1 X8Y0VDDM 20mOhm
LX8Y0VDD X8Y0VDDM VDD2 0.036nH
RX8Y0VSS VSS1 X8Y0VSSM 20mOhm
LX8Y0VSS X8Y0VSSM VSS2 0.036nH
RX8Y1VDD VDD1 X8Y1VDDM 20mOhm
LX8Y1VDD X8Y1VDDM VDD2 0.036nH
RX8Y1VSS VSS1 X8Y1VSSM 20mOhm
LX8Y1VSS X8Y1VSSM VSS2 0.036nH
RX8Y2VDD VDD1 X8Y2VDDM 20mOhm
LX8Y2VDD X8Y2VDDM VDD2 0.036nH
RX8Y2VSS VSS1 X8Y2VSSM 20mOhm
LX8Y2VSS X8Y2VSSM VSS2 0.036nH
RX8Y3VDD VDD1 X8Y3VDDM 20mOhm
LX8Y3VDD X8Y3VDDM VDD2 0.036nH
RX8Y3VSS VSS1 X8Y3VSSM 20mOhm
LX8Y3VSS X8Y3VSSM VSS2 0.036nH
RX8Y4VDD VDD1 X8Y4VDDM 20mOhm
LX8Y4VDD X8Y4VDDM VDD2 0.036nH
RX8Y4VSS VSS1 X8Y4VSSM 20mOhm
LX8Y4VSS X8Y4VSSM VSS2 0.036nH
RX8Y5VDD VDD1 X8Y5VDDM 20mOhm
LX8Y5VDD X8Y5VDDM VDD2 0.036nH
RX8Y5VSS VSS1 X8Y5VSSM 20mOhm
LX8Y5VSS X8Y5VSSM VSS2 0.036nH
RX8Y6VDD VDD1 X8Y6VDDM 20mOhm
LX8Y6VDD X8Y6VDDM VDD2 0.036nH
RX8Y6VSS VSS1 X8Y6VSSM 20mOhm
LX8Y6VSS X8Y6VSSM VSS2 0.036nH
RX8Y7VDD VDD1 X8Y7VDDM 20mOhm
LX8Y7VDD X8Y7VDDM VDD2 0.036nH
RX8Y7VSS VSS1 X8Y7VSSM 20mOhm
LX8Y7VSS X8Y7VSSM VSS2 0.036nH
RX8Y8VDD VDD1 X8Y8VDDM 20mOhm
LX8Y8VDD X8Y8VDDM VDD2 0.036nH
RX8Y8VSS VSS1 X8Y8VSSM 20mOhm
LX8Y8VSS X8Y8VSSM VSS2 0.036nH
RX8Y9VDD VDD1 X8Y9VDDM 20mOhm
LX8Y9VDD X8Y9VDDM VDD2 0.036nH
RX8Y9VSS VSS1 X8Y9VSSM 20mOhm
LX8Y9VSS X8Y9VSSM VSS2 0.036nH
RX8Y10VDD VDD1 X8Y10VDDM 20mOhm
LX8Y10VDD X8Y10VDDM VDD2 0.036nH
RX8Y10VSS VSS1 X8Y10VSSM 20mOhm
LX8Y10VSS X8Y10VSSM VSS2 0.036nH
RX8Y11VDD VDD1 X8Y11VDDM 20mOhm
LX8Y11VDD X8Y11VDDM VDD2 0.036nH
RX8Y11VSS VSS1 X8Y11VSSM 20mOhm
LX8Y11VSS X8Y11VSSM VSS2 0.036nH
RX9Y0VDD VDD1 X9Y0VDDM 20mOhm
LX9Y0VDD X9Y0VDDM VDD2 0.036nH
RX9Y0VSS VSS1 X9Y0VSSM 20mOhm
LX9Y0VSS X9Y0VSSM VSS2 0.036nH
RX9Y1VDD VDD1 X9Y1VDDM 20mOhm
LX9Y1VDD X9Y1VDDM VDD2 0.036nH
RX9Y1VSS VSS1 X9Y1VSSM 20mOhm
LX9Y1VSS X9Y1VSSM VSS2 0.036nH
RX9Y2VDD VDD1 X9Y2VDDM 20mOhm
LX9Y2VDD X9Y2VDDM VDD2 0.036nH
RX9Y2VSS VSS1 X9Y2VSSM 20mOhm
LX9Y2VSS X9Y2VSSM VSS2 0.036nH
RX9Y3VDD VDD1 X9Y3VDDM 20mOhm
LX9Y3VDD X9Y3VDDM VDD2 0.036nH
RX9Y3VSS VSS1 X9Y3VSSM 20mOhm
LX9Y3VSS X9Y3VSSM VSS2 0.036nH
RX9Y4VDD VDD1 X9Y4VDDM 20mOhm
LX9Y4VDD X9Y4VDDM VDD2 0.036nH
RX9Y4VSS VSS1 X9Y4VSSM 20mOhm
LX9Y4VSS X9Y4VSSM VSS2 0.036nH
RX9Y5VDD VDD1 X9Y5VDDM 20mOhm
LX9Y5VDD X9Y5VDDM VDD2 0.036nH
RX9Y5VSS VSS1 X9Y5VSSM 20mOhm
LX9Y5VSS X9Y5VSSM VSS2 0.036nH
RX9Y6VDD VDD1 X9Y6VDDM 20mOhm
LX9Y6VDD X9Y6VDDM VDD2 0.036nH
RX9Y6VSS VSS1 X9Y6VSSM 20mOhm
LX9Y6VSS X9Y6VSSM VSS2 0.036nH
RX9Y7VDD VDD1 X9Y7VDDM 20mOhm
LX9Y7VDD X9Y7VDDM VDD2 0.036nH
RX9Y7VSS VSS1 X9Y7VSSM 20mOhm
LX9Y7VSS X9Y7VSSM VSS2 0.036nH
RX9Y8VDD VDD1 X9Y8VDDM 20mOhm
LX9Y8VDD X9Y8VDDM VDD2 0.036nH
RX9Y8VSS VSS1 X9Y8VSSM 20mOhm
LX9Y8VSS X9Y8VSSM VSS2 0.036nH
RX9Y9VDD VDD1 X9Y9VDDM 20mOhm
LX9Y9VDD X9Y9VDDM VDD2 0.036nH
RX9Y9VSS VSS1 X9Y9VSSM 20mOhm
LX9Y9VSS X9Y9VSSM VSS2 0.036nH
RX9Y10VDD VDD1 X9Y10VDDM 20mOhm
LX9Y10VDD X9Y10VDDM VDD2 0.036nH
RX9Y10VSS VSS1 X9Y10VSSM 20mOhm
LX9Y10VSS X9Y10VSSM VSS2 0.036nH
RX9Y11VDD VDD1 X9Y11VDDM 20mOhm
LX9Y11VDD X9Y11VDDM VDD2 0.036nH
RX9Y11VSS VSS1 X9Y11VSSM 20mOhm
LX9Y11VSS X9Y11VSSM VSS2 0.036nH
RX10Y0VDD VDD1 X10Y0VDDM 20mOhm
LX10Y0VDD X10Y0VDDM VDD2 0.036nH
RX10Y0VSS VSS1 X10Y0VSSM 20mOhm
LX10Y0VSS X10Y0VSSM VSS2 0.036nH
RX10Y1VDD VDD1 X10Y1VDDM 20mOhm
LX10Y1VDD X10Y1VDDM VDD2 0.036nH
RX10Y1VSS VSS1 X10Y1VSSM 20mOhm
LX10Y1VSS X10Y1VSSM VSS2 0.036nH
RX10Y2VDD VDD1 X10Y2VDDM 20mOhm
LX10Y2VDD X10Y2VDDM VDD2 0.036nH
RX10Y2VSS VSS1 X10Y2VSSM 20mOhm
LX10Y2VSS X10Y2VSSM VSS2 0.036nH
RX10Y3VDD VDD1 X10Y3VDDM 20mOhm
LX10Y3VDD X10Y3VDDM VDD2 0.036nH
RX10Y3VSS VSS1 X10Y3VSSM 20mOhm
LX10Y3VSS X10Y3VSSM VSS2 0.036nH
RX10Y4VDD VDD1 X10Y4VDDM 20mOhm
LX10Y4VDD X10Y4VDDM VDD2 0.036nH
RX10Y4VSS VSS1 X10Y4VSSM 20mOhm
LX10Y4VSS X10Y4VSSM VSS2 0.036nH
RX10Y5VDD VDD1 X10Y5VDDM 20mOhm
LX10Y5VDD X10Y5VDDM VDD2 0.036nH
RX10Y5VSS VSS1 X10Y5VSSM 20mOhm
LX10Y5VSS X10Y5VSSM VSS2 0.036nH
RX10Y6VDD VDD1 X10Y6VDDM 20mOhm
LX10Y6VDD X10Y6VDDM VDD2 0.036nH
RX10Y6VSS VSS1 X10Y6VSSM 20mOhm
LX10Y6VSS X10Y6VSSM VSS2 0.036nH
RX10Y7VDD VDD1 X10Y7VDDM 20mOhm
LX10Y7VDD X10Y7VDDM VDD2 0.036nH
RX10Y7VSS VSS1 X10Y7VSSM 20mOhm
LX10Y7VSS X10Y7VSSM VSS2 0.036nH
RX10Y8VDD VDD1 X10Y8VDDM 20mOhm
LX10Y8VDD X10Y8VDDM VDD2 0.036nH
RX10Y8VSS VSS1 X10Y8VSSM 20mOhm
LX10Y8VSS X10Y8VSSM VSS2 0.036nH
RX10Y9VDD VDD1 X10Y9VDDM 20mOhm
LX10Y9VDD X10Y9VDDM VDD2 0.036nH
RX10Y9VSS VSS1 X10Y9VSSM 20mOhm
LX10Y9VSS X10Y9VSSM VSS2 0.036nH
RX10Y10VDD VDD1 X10Y10VDDM 20mOhm
LX10Y10VDD X10Y10VDDM VDD2 0.036nH
RX10Y10VSS VSS1 X10Y10VSSM 20mOhm
LX10Y10VSS X10Y10VSSM VSS2 0.036nH
RX10Y11VDD VDD1 X10Y11VDDM 20mOhm
LX10Y11VDD X10Y11VDDM VDD2 0.036nH
RX10Y11VSS VSS1 X10Y11VSSM 20mOhm
LX10Y11VSS X10Y11VSSM VSS2 0.036nH
RX11Y0VDD VDD1 X11Y0VDDM 20mOhm
LX11Y0VDD X11Y0VDDM VDD2 0.036nH
RX11Y0VSS VSS1 X11Y0VSSM 20mOhm
LX11Y0VSS X11Y0VSSM VSS2 0.036nH
RX11Y1VDD VDD1 X11Y1VDDM 20mOhm
LX11Y1VDD X11Y1VDDM VDD2 0.036nH
RX11Y1VSS VSS1 X11Y1VSSM 20mOhm
LX11Y1VSS X11Y1VSSM VSS2 0.036nH
RX11Y2VDD VDD1 X11Y2VDDM 20mOhm
LX11Y2VDD X11Y2VDDM VDD2 0.036nH
RX11Y2VSS VSS1 X11Y2VSSM 20mOhm
LX11Y2VSS X11Y2VSSM VSS2 0.036nH
RX11Y3VDD VDD1 X11Y3VDDM 20mOhm
LX11Y3VDD X11Y3VDDM VDD2 0.036nH
RX11Y3VSS VSS1 X11Y3VSSM 20mOhm
LX11Y3VSS X11Y3VSSM VSS2 0.036nH
RX11Y4VDD VDD1 X11Y4VDDM 20mOhm
LX11Y4VDD X11Y4VDDM VDD2 0.036nH
RX11Y4VSS VSS1 X11Y4VSSM 20mOhm
LX11Y4VSS X11Y4VSSM VSS2 0.036nH
RX11Y5VDD VDD1 X11Y5VDDM 20mOhm
LX11Y5VDD X11Y5VDDM VDD2 0.036nH
RX11Y5VSS VSS1 X11Y5VSSM 20mOhm
LX11Y5VSS X11Y5VSSM VSS2 0.036nH
RX11Y6VDD VDD1 X11Y6VDDM 20mOhm
LX11Y6VDD X11Y6VDDM VDD2 0.036nH
RX11Y6VSS VSS1 X11Y6VSSM 20mOhm
LX11Y6VSS X11Y6VSSM VSS2 0.036nH
RX11Y7VDD VDD1 X11Y7VDDM 20mOhm
LX11Y7VDD X11Y7VDDM VDD2 0.036nH
RX11Y7VSS VSS1 X11Y7VSSM 20mOhm
LX11Y7VSS X11Y7VSSM VSS2 0.036nH
RX11Y8VDD VDD1 X11Y8VDDM 20mOhm
LX11Y8VDD X11Y8VDDM VDD2 0.036nH
RX11Y8VSS VSS1 X11Y8VSSM 20mOhm
LX11Y8VSS X11Y8VSSM VSS2 0.036nH
RX11Y9VDD VDD1 X11Y9VDDM 20mOhm
LX11Y9VDD X11Y9VDDM VDD2 0.036nH
RX11Y9VSS VSS1 X11Y9VSSM 20mOhm
LX11Y9VSS X11Y9VSSM VSS2 0.036nH
RX11Y10VDD VDD1 X11Y10VDDM 20mOhm
LX11Y10VDD X11Y10VDDM VDD2 0.036nH
RX11Y10VSS VSS1 X11Y10VSSM 20mOhm
LX11Y10VSS X11Y10VSSM VSS2 0.036nH
RX11Y11VDD VDD1 X11Y11VDDM 20mOhm
LX11Y11VDD X11Y11VDDM VDD2 0.036nH
RX11Y11VSS VSS1 X11Y11VSSM 20mOhm
LX11Y11VSS X11Y11VSSM VSS2 0.036nH
.ends ChipBump

.subckt PcbModelLumped VDD1 VSS1 VDD2 VSS2
Rs1 VDD1 11 1000mOhm
Ls1 11 VDD2 0nH
Rs2 VSS1 21 1000mOhm
Ls2 21 VSS2 0nH
Rp VDD2 VDD2M 0mOhm
Cp VDD2M VSS2 0uF
.ends PcbModelLumped

.subckt dut VDD VSS
R_X10Y10VDD_X20Y10VDD X10Y10VDD X15Y10VDD 25mOhm
L_X10Y10VDD_X20Y10VDD X15Y10VDD X20Y10VDD 2.91e-06nH
R_X10Y10VSS_X20Y10VSS X10Y10VSS X15Y10VSS 25mOhm
L_X10Y10VSS_X20Y10VSS X15Y10VSS X20Y10VSS 2.91e-06nH
R_X20Y10VDD_X30Y10VDD X20Y10VDD X25Y10VDD 25mOhm
L_X20Y10VDD_X30Y10VDD X25Y10VDD X30Y10VDD 2.91e-06nH
R_X20Y10VSS_X30Y10VSS X20Y10VSS X25Y10VSS 25mOhm
L_X20Y10VSS_X30Y10VSS X25Y10VSS X30Y10VSS 2.91e-06nH
R_X30Y10VDD_X40Y10VDD X30Y10VDD X35Y10VDD 25mOhm
L_X30Y10VDD_X40Y10VDD X35Y10VDD X40Y10VDD 2.91e-06nH
R_X30Y10VSS_X40Y10VSS X30Y10VSS X35Y10VSS 25mOhm
L_X30Y10VSS_X40Y10VSS X35Y10VSS X40Y10VSS 2.91e-06nH
R_X40Y10VDD_X50Y10VDD X40Y10VDD X45Y10VDD 25mOhm
L_X40Y10VDD_X50Y10VDD X45Y10VDD X50Y10VDD 2.91e-06nH
R_X40Y10VSS_X50Y10VSS X40Y10VSS X45Y10VSS 25mOhm
L_X40Y10VSS_X50Y10VSS X45Y10VSS X50Y10VSS 2.91e-06nH
R_X50Y10VDD_X60Y10VDD X50Y10VDD X55Y10VDD 25mOhm
L_X50Y10VDD_X60Y10VDD X55Y10VDD X60Y10VDD 2.91e-06nH
R_X50Y10VSS_X60Y10VSS X50Y10VSS X55Y10VSS 25mOhm
L_X50Y10VSS_X60Y10VSS X55Y10VSS X60Y10VSS 2.91e-06nH
R_X60Y10VDD_X70Y10VDD X60Y10VDD X65Y10VDD 25mOhm
L_X60Y10VDD_X70Y10VDD X65Y10VDD X70Y10VDD 2.91e-06nH
R_X60Y10VSS_X70Y10VSS X60Y10VSS X65Y10VSS 25mOhm
L_X60Y10VSS_X70Y10VSS X65Y10VSS X70Y10VSS 2.91e-06nH
R_X70Y10VDD_X80Y10VDD X70Y10VDD X75Y10VDD 25mOhm
L_X70Y10VDD_X80Y10VDD X75Y10VDD X80Y10VDD 2.91e-06nH
R_X70Y10VSS_X80Y10VSS X70Y10VSS X75Y10VSS 25mOhm
L_X70Y10VSS_X80Y10VSS X75Y10VSS X80Y10VSS 2.91e-06nH
R_X80Y10VDD_X90Y10VDD X80Y10VDD X85Y10VDD 25mOhm
L_X80Y10VDD_X90Y10VDD X85Y10VDD X90Y10VDD 2.91e-06nH
R_X80Y10VSS_X90Y10VSS X80Y10VSS X85Y10VSS 25mOhm
L_X80Y10VSS_X90Y10VSS X85Y10VSS X90Y10VSS 2.91e-06nH
R_X90Y10VDD_X100Y10VDD X90Y10VDD X95Y10VDD 25mOhm
L_X90Y10VDD_X100Y10VDD X95Y10VDD X100Y10VDD 2.91e-06nH
R_X90Y10VSS_X100Y10VSS X90Y10VSS X95Y10VSS 25mOhm
L_X90Y10VSS_X100Y10VSS X95Y10VSS X100Y10VSS 2.91e-06nH
R_X100Y10VDD_X110Y10VDD X100Y10VDD X105Y10VDD 25mOhm
L_X100Y10VDD_X110Y10VDD X105Y10VDD X110Y10VDD 2.91e-06nH
R_X100Y10VSS_X110Y10VSS X100Y10VSS X105Y10VSS 25mOhm
L_X100Y10VSS_X110Y10VSS X105Y10VSS X110Y10VSS 2.91e-06nH
R_X110Y10VDD_X120Y10VDD X110Y10VDD X115Y10VDD 25mOhm
L_X110Y10VDD_X120Y10VDD X115Y10VDD X120Y10VDD 2.91e-06nH
R_X110Y10VSS_X120Y10VSS X110Y10VSS X115Y10VSS 25mOhm
L_X110Y10VSS_X120Y10VSS X115Y10VSS X120Y10VSS 2.91e-06nH
R_X10Y20VDD_X20Y20VDD X10Y20VDD X15Y20VDD 25mOhm
L_X10Y20VDD_X20Y20VDD X15Y20VDD X20Y20VDD 2.91e-06nH
R_X10Y20VSS_X20Y20VSS X10Y20VSS X15Y20VSS 25mOhm
L_X10Y20VSS_X20Y20VSS X15Y20VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X30Y20VDD X20Y20VDD X25Y20VDD 25mOhm
L_X20Y20VDD_X30Y20VDD X25Y20VDD X30Y20VDD 2.91e-06nH
R_X20Y20VSS_X30Y20VSS X20Y20VSS X25Y20VSS 25mOhm
L_X20Y20VSS_X30Y20VSS X25Y20VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X40Y20VDD X30Y20VDD X35Y20VDD 25mOhm
L_X30Y20VDD_X40Y20VDD X35Y20VDD X40Y20VDD 2.91e-06nH
R_X30Y20VSS_X40Y20VSS X30Y20VSS X35Y20VSS 25mOhm
L_X30Y20VSS_X40Y20VSS X35Y20VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X50Y20VDD X40Y20VDD X45Y20VDD 25mOhm
L_X40Y20VDD_X50Y20VDD X45Y20VDD X50Y20VDD 2.91e-06nH
R_X40Y20VSS_X50Y20VSS X40Y20VSS X45Y20VSS 25mOhm
L_X40Y20VSS_X50Y20VSS X45Y20VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X60Y20VDD X50Y20VDD X55Y20VDD 25mOhm
L_X50Y20VDD_X60Y20VDD X55Y20VDD X60Y20VDD 2.91e-06nH
R_X50Y20VSS_X60Y20VSS X50Y20VSS X55Y20VSS 25mOhm
L_X50Y20VSS_X60Y20VSS X55Y20VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X70Y20VDD X60Y20VDD X65Y20VDD 25mOhm
L_X60Y20VDD_X70Y20VDD X65Y20VDD X70Y20VDD 2.91e-06nH
R_X60Y20VSS_X70Y20VSS X60Y20VSS X65Y20VSS 25mOhm
L_X60Y20VSS_X70Y20VSS X65Y20VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X80Y20VDD X70Y20VDD X75Y20VDD 25mOhm
L_X70Y20VDD_X80Y20VDD X75Y20VDD X80Y20VDD 2.91e-06nH
R_X70Y20VSS_X80Y20VSS X70Y20VSS X75Y20VSS 25mOhm
L_X70Y20VSS_X80Y20VSS X75Y20VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X90Y20VDD X80Y20VDD X85Y20VDD 25mOhm
L_X80Y20VDD_X90Y20VDD X85Y20VDD X90Y20VDD 2.91e-06nH
R_X80Y20VSS_X90Y20VSS X80Y20VSS X85Y20VSS 25mOhm
L_X80Y20VSS_X90Y20VSS X85Y20VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X100Y20VDD X90Y20VDD X95Y20VDD 25mOhm
L_X90Y20VDD_X100Y20VDD X95Y20VDD X100Y20VDD 2.91e-06nH
R_X90Y20VSS_X100Y20VSS X90Y20VSS X95Y20VSS 25mOhm
L_X90Y20VSS_X100Y20VSS X95Y20VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X110Y20VDD X100Y20VDD X105Y20VDD 25mOhm
L_X100Y20VDD_X110Y20VDD X105Y20VDD X110Y20VDD 2.91e-06nH
R_X100Y20VSS_X110Y20VSS X100Y20VSS X105Y20VSS 25mOhm
L_X100Y20VSS_X110Y20VSS X105Y20VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X120Y20VDD X110Y20VDD X115Y20VDD 25mOhm
L_X110Y20VDD_X120Y20VDD X115Y20VDD X120Y20VDD 2.91e-06nH
R_X110Y20VSS_X120Y20VSS X110Y20VSS X115Y20VSS 25mOhm
L_X110Y20VSS_X120Y20VSS X115Y20VSS X120Y20VSS 2.91e-06nH
R_X10Y30VDD_X20Y30VDD X10Y30VDD X15Y30VDD 25mOhm
L_X10Y30VDD_X20Y30VDD X15Y30VDD X20Y30VDD 2.91e-06nH
R_X10Y30VSS_X20Y30VSS X10Y30VSS X15Y30VSS 25mOhm
L_X10Y30VSS_X20Y30VSS X15Y30VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X30Y30VDD X20Y30VDD X25Y30VDD 25mOhm
L_X20Y30VDD_X30Y30VDD X25Y30VDD X30Y30VDD 2.91e-06nH
R_X20Y30VSS_X30Y30VSS X20Y30VSS X25Y30VSS 25mOhm
L_X20Y30VSS_X30Y30VSS X25Y30VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X40Y30VDD X30Y30VDD X35Y30VDD 25mOhm
L_X30Y30VDD_X40Y30VDD X35Y30VDD X40Y30VDD 2.91e-06nH
R_X30Y30VSS_X40Y30VSS X30Y30VSS X35Y30VSS 25mOhm
L_X30Y30VSS_X40Y30VSS X35Y30VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X50Y30VDD X40Y30VDD X45Y30VDD 25mOhm
L_X40Y30VDD_X50Y30VDD X45Y30VDD X50Y30VDD 2.91e-06nH
R_X40Y30VSS_X50Y30VSS X40Y30VSS X45Y30VSS 25mOhm
L_X40Y30VSS_X50Y30VSS X45Y30VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X60Y30VDD X50Y30VDD X55Y30VDD 25mOhm
L_X50Y30VDD_X60Y30VDD X55Y30VDD X60Y30VDD 2.91e-06nH
R_X50Y30VSS_X60Y30VSS X50Y30VSS X55Y30VSS 25mOhm
L_X50Y30VSS_X60Y30VSS X55Y30VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X70Y30VDD X60Y30VDD X65Y30VDD 25mOhm
L_X60Y30VDD_X70Y30VDD X65Y30VDD X70Y30VDD 2.91e-06nH
R_X60Y30VSS_X70Y30VSS X60Y30VSS X65Y30VSS 25mOhm
L_X60Y30VSS_X70Y30VSS X65Y30VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X80Y30VDD X70Y30VDD X75Y30VDD 25mOhm
L_X70Y30VDD_X80Y30VDD X75Y30VDD X80Y30VDD 2.91e-06nH
R_X70Y30VSS_X80Y30VSS X70Y30VSS X75Y30VSS 25mOhm
L_X70Y30VSS_X80Y30VSS X75Y30VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X90Y30VDD X80Y30VDD X85Y30VDD 25mOhm
L_X80Y30VDD_X90Y30VDD X85Y30VDD X90Y30VDD 2.91e-06nH
R_X80Y30VSS_X90Y30VSS X80Y30VSS X85Y30VSS 25mOhm
L_X80Y30VSS_X90Y30VSS X85Y30VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X100Y30VDD X90Y30VDD X95Y30VDD 25mOhm
L_X90Y30VDD_X100Y30VDD X95Y30VDD X100Y30VDD 2.91e-06nH
R_X90Y30VSS_X100Y30VSS X90Y30VSS X95Y30VSS 25mOhm
L_X90Y30VSS_X100Y30VSS X95Y30VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X110Y30VDD X100Y30VDD X105Y30VDD 25mOhm
L_X100Y30VDD_X110Y30VDD X105Y30VDD X110Y30VDD 2.91e-06nH
R_X100Y30VSS_X110Y30VSS X100Y30VSS X105Y30VSS 25mOhm
L_X100Y30VSS_X110Y30VSS X105Y30VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X120Y30VDD X110Y30VDD X115Y30VDD 25mOhm
L_X110Y30VDD_X120Y30VDD X115Y30VDD X120Y30VDD 2.91e-06nH
R_X110Y30VSS_X120Y30VSS X110Y30VSS X115Y30VSS 25mOhm
L_X110Y30VSS_X120Y30VSS X115Y30VSS X120Y30VSS 2.91e-06nH
R_X10Y40VDD_X20Y40VDD X10Y40VDD X15Y40VDD 25mOhm
L_X10Y40VDD_X20Y40VDD X15Y40VDD X20Y40VDD 2.91e-06nH
R_X10Y40VSS_X20Y40VSS X10Y40VSS X15Y40VSS 25mOhm
L_X10Y40VSS_X20Y40VSS X15Y40VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X30Y40VDD X20Y40VDD X25Y40VDD 25mOhm
L_X20Y40VDD_X30Y40VDD X25Y40VDD X30Y40VDD 2.91e-06nH
R_X20Y40VSS_X30Y40VSS X20Y40VSS X25Y40VSS 25mOhm
L_X20Y40VSS_X30Y40VSS X25Y40VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X40Y40VDD X30Y40VDD X35Y40VDD 25mOhm
L_X30Y40VDD_X40Y40VDD X35Y40VDD X40Y40VDD 2.91e-06nH
R_X30Y40VSS_X40Y40VSS X30Y40VSS X35Y40VSS 25mOhm
L_X30Y40VSS_X40Y40VSS X35Y40VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X50Y40VDD X40Y40VDD X45Y40VDD 25mOhm
L_X40Y40VDD_X50Y40VDD X45Y40VDD X50Y40VDD 2.91e-06nH
R_X40Y40VSS_X50Y40VSS X40Y40VSS X45Y40VSS 25mOhm
L_X40Y40VSS_X50Y40VSS X45Y40VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X60Y40VDD X50Y40VDD X55Y40VDD 25mOhm
L_X50Y40VDD_X60Y40VDD X55Y40VDD X60Y40VDD 2.91e-06nH
R_X50Y40VSS_X60Y40VSS X50Y40VSS X55Y40VSS 25mOhm
L_X50Y40VSS_X60Y40VSS X55Y40VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X70Y40VDD X60Y40VDD X65Y40VDD 25mOhm
L_X60Y40VDD_X70Y40VDD X65Y40VDD X70Y40VDD 2.91e-06nH
R_X60Y40VSS_X70Y40VSS X60Y40VSS X65Y40VSS 25mOhm
L_X60Y40VSS_X70Y40VSS X65Y40VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X80Y40VDD X70Y40VDD X75Y40VDD 25mOhm
L_X70Y40VDD_X80Y40VDD X75Y40VDD X80Y40VDD 2.91e-06nH
R_X70Y40VSS_X80Y40VSS X70Y40VSS X75Y40VSS 25mOhm
L_X70Y40VSS_X80Y40VSS X75Y40VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X90Y40VDD X80Y40VDD X85Y40VDD 25mOhm
L_X80Y40VDD_X90Y40VDD X85Y40VDD X90Y40VDD 2.91e-06nH
R_X80Y40VSS_X90Y40VSS X80Y40VSS X85Y40VSS 25mOhm
L_X80Y40VSS_X90Y40VSS X85Y40VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X100Y40VDD X90Y40VDD X95Y40VDD 25mOhm
L_X90Y40VDD_X100Y40VDD X95Y40VDD X100Y40VDD 2.91e-06nH
R_X90Y40VSS_X100Y40VSS X90Y40VSS X95Y40VSS 25mOhm
L_X90Y40VSS_X100Y40VSS X95Y40VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X110Y40VDD X100Y40VDD X105Y40VDD 25mOhm
L_X100Y40VDD_X110Y40VDD X105Y40VDD X110Y40VDD 2.91e-06nH
R_X100Y40VSS_X110Y40VSS X100Y40VSS X105Y40VSS 25mOhm
L_X100Y40VSS_X110Y40VSS X105Y40VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X120Y40VDD X110Y40VDD X115Y40VDD 25mOhm
L_X110Y40VDD_X120Y40VDD X115Y40VDD X120Y40VDD 2.91e-06nH
R_X110Y40VSS_X120Y40VSS X110Y40VSS X115Y40VSS 25mOhm
L_X110Y40VSS_X120Y40VSS X115Y40VSS X120Y40VSS 2.91e-06nH
R_X10Y50VDD_X20Y50VDD X10Y50VDD X15Y50VDD 25mOhm
L_X10Y50VDD_X20Y50VDD X15Y50VDD X20Y50VDD 2.91e-06nH
R_X10Y50VSS_X20Y50VSS X10Y50VSS X15Y50VSS 25mOhm
L_X10Y50VSS_X20Y50VSS X15Y50VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X30Y50VDD X20Y50VDD X25Y50VDD 25mOhm
L_X20Y50VDD_X30Y50VDD X25Y50VDD X30Y50VDD 2.91e-06nH
R_X20Y50VSS_X30Y50VSS X20Y50VSS X25Y50VSS 25mOhm
L_X20Y50VSS_X30Y50VSS X25Y50VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X40Y50VDD X30Y50VDD X35Y50VDD 25mOhm
L_X30Y50VDD_X40Y50VDD X35Y50VDD X40Y50VDD 2.91e-06nH
R_X30Y50VSS_X40Y50VSS X30Y50VSS X35Y50VSS 25mOhm
L_X30Y50VSS_X40Y50VSS X35Y50VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X50Y50VDD X40Y50VDD X45Y50VDD 25mOhm
L_X40Y50VDD_X50Y50VDD X45Y50VDD X50Y50VDD 2.91e-06nH
R_X40Y50VSS_X50Y50VSS X40Y50VSS X45Y50VSS 25mOhm
L_X40Y50VSS_X50Y50VSS X45Y50VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X60Y50VDD X50Y50VDD X55Y50VDD 25mOhm
L_X50Y50VDD_X60Y50VDD X55Y50VDD X60Y50VDD 2.91e-06nH
R_X50Y50VSS_X60Y50VSS X50Y50VSS X55Y50VSS 25mOhm
L_X50Y50VSS_X60Y50VSS X55Y50VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X70Y50VDD X60Y50VDD X65Y50VDD 25mOhm
L_X60Y50VDD_X70Y50VDD X65Y50VDD X70Y50VDD 2.91e-06nH
R_X60Y50VSS_X70Y50VSS X60Y50VSS X65Y50VSS 25mOhm
L_X60Y50VSS_X70Y50VSS X65Y50VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X80Y50VDD X70Y50VDD X75Y50VDD 25mOhm
L_X70Y50VDD_X80Y50VDD X75Y50VDD X80Y50VDD 2.91e-06nH
R_X70Y50VSS_X80Y50VSS X70Y50VSS X75Y50VSS 25mOhm
L_X70Y50VSS_X80Y50VSS X75Y50VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X90Y50VDD X80Y50VDD X85Y50VDD 25mOhm
L_X80Y50VDD_X90Y50VDD X85Y50VDD X90Y50VDD 2.91e-06nH
R_X80Y50VSS_X90Y50VSS X80Y50VSS X85Y50VSS 25mOhm
L_X80Y50VSS_X90Y50VSS X85Y50VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X100Y50VDD X90Y50VDD X95Y50VDD 25mOhm
L_X90Y50VDD_X100Y50VDD X95Y50VDD X100Y50VDD 2.91e-06nH
R_X90Y50VSS_X100Y50VSS X90Y50VSS X95Y50VSS 25mOhm
L_X90Y50VSS_X100Y50VSS X95Y50VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X110Y50VDD X100Y50VDD X105Y50VDD 25mOhm
L_X100Y50VDD_X110Y50VDD X105Y50VDD X110Y50VDD 2.91e-06nH
R_X100Y50VSS_X110Y50VSS X100Y50VSS X105Y50VSS 25mOhm
L_X100Y50VSS_X110Y50VSS X105Y50VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X120Y50VDD X110Y50VDD X115Y50VDD 25mOhm
L_X110Y50VDD_X120Y50VDD X115Y50VDD X120Y50VDD 2.91e-06nH
R_X110Y50VSS_X120Y50VSS X110Y50VSS X115Y50VSS 25mOhm
L_X110Y50VSS_X120Y50VSS X115Y50VSS X120Y50VSS 2.91e-06nH
R_X10Y60VDD_X20Y60VDD X10Y60VDD X15Y60VDD 25mOhm
L_X10Y60VDD_X20Y60VDD X15Y60VDD X20Y60VDD 2.91e-06nH
R_X10Y60VSS_X20Y60VSS X10Y60VSS X15Y60VSS 25mOhm
L_X10Y60VSS_X20Y60VSS X15Y60VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X30Y60VDD X20Y60VDD X25Y60VDD 25mOhm
L_X20Y60VDD_X30Y60VDD X25Y60VDD X30Y60VDD 2.91e-06nH
R_X20Y60VSS_X30Y60VSS X20Y60VSS X25Y60VSS 25mOhm
L_X20Y60VSS_X30Y60VSS X25Y60VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X40Y60VDD X30Y60VDD X35Y60VDD 25mOhm
L_X30Y60VDD_X40Y60VDD X35Y60VDD X40Y60VDD 2.91e-06nH
R_X30Y60VSS_X40Y60VSS X30Y60VSS X35Y60VSS 25mOhm
L_X30Y60VSS_X40Y60VSS X35Y60VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X50Y60VDD X40Y60VDD X45Y60VDD 25mOhm
L_X40Y60VDD_X50Y60VDD X45Y60VDD X50Y60VDD 2.91e-06nH
R_X40Y60VSS_X50Y60VSS X40Y60VSS X45Y60VSS 25mOhm
L_X40Y60VSS_X50Y60VSS X45Y60VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X60Y60VDD X50Y60VDD X55Y60VDD 25mOhm
L_X50Y60VDD_X60Y60VDD X55Y60VDD X60Y60VDD 2.91e-06nH
R_X50Y60VSS_X60Y60VSS X50Y60VSS X55Y60VSS 25mOhm
L_X50Y60VSS_X60Y60VSS X55Y60VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X70Y60VDD X60Y60VDD X65Y60VDD 25mOhm
L_X60Y60VDD_X70Y60VDD X65Y60VDD X70Y60VDD 2.91e-06nH
R_X60Y60VSS_X70Y60VSS X60Y60VSS X65Y60VSS 25mOhm
L_X60Y60VSS_X70Y60VSS X65Y60VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X80Y60VDD X70Y60VDD X75Y60VDD 25mOhm
L_X70Y60VDD_X80Y60VDD X75Y60VDD X80Y60VDD 2.91e-06nH
R_X70Y60VSS_X80Y60VSS X70Y60VSS X75Y60VSS 25mOhm
L_X70Y60VSS_X80Y60VSS X75Y60VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X90Y60VDD X80Y60VDD X85Y60VDD 25mOhm
L_X80Y60VDD_X90Y60VDD X85Y60VDD X90Y60VDD 2.91e-06nH
R_X80Y60VSS_X90Y60VSS X80Y60VSS X85Y60VSS 25mOhm
L_X80Y60VSS_X90Y60VSS X85Y60VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X100Y60VDD X90Y60VDD X95Y60VDD 25mOhm
L_X90Y60VDD_X100Y60VDD X95Y60VDD X100Y60VDD 2.91e-06nH
R_X90Y60VSS_X100Y60VSS X90Y60VSS X95Y60VSS 25mOhm
L_X90Y60VSS_X100Y60VSS X95Y60VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X110Y60VDD X100Y60VDD X105Y60VDD 25mOhm
L_X100Y60VDD_X110Y60VDD X105Y60VDD X110Y60VDD 2.91e-06nH
R_X100Y60VSS_X110Y60VSS X100Y60VSS X105Y60VSS 25mOhm
L_X100Y60VSS_X110Y60VSS X105Y60VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X120Y60VDD X110Y60VDD X115Y60VDD 25mOhm
L_X110Y60VDD_X120Y60VDD X115Y60VDD X120Y60VDD 2.91e-06nH
R_X110Y60VSS_X120Y60VSS X110Y60VSS X115Y60VSS 25mOhm
L_X110Y60VSS_X120Y60VSS X115Y60VSS X120Y60VSS 2.91e-06nH
R_X10Y70VDD_X20Y70VDD X10Y70VDD X15Y70VDD 25mOhm
L_X10Y70VDD_X20Y70VDD X15Y70VDD X20Y70VDD 2.91e-06nH
R_X10Y70VSS_X20Y70VSS X10Y70VSS X15Y70VSS 25mOhm
L_X10Y70VSS_X20Y70VSS X15Y70VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X30Y70VDD X20Y70VDD X25Y70VDD 25mOhm
L_X20Y70VDD_X30Y70VDD X25Y70VDD X30Y70VDD 2.91e-06nH
R_X20Y70VSS_X30Y70VSS X20Y70VSS X25Y70VSS 25mOhm
L_X20Y70VSS_X30Y70VSS X25Y70VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X40Y70VDD X30Y70VDD X35Y70VDD 25mOhm
L_X30Y70VDD_X40Y70VDD X35Y70VDD X40Y70VDD 2.91e-06nH
R_X30Y70VSS_X40Y70VSS X30Y70VSS X35Y70VSS 25mOhm
L_X30Y70VSS_X40Y70VSS X35Y70VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X50Y70VDD X40Y70VDD X45Y70VDD 25mOhm
L_X40Y70VDD_X50Y70VDD X45Y70VDD X50Y70VDD 2.91e-06nH
R_X40Y70VSS_X50Y70VSS X40Y70VSS X45Y70VSS 25mOhm
L_X40Y70VSS_X50Y70VSS X45Y70VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X60Y70VDD X50Y70VDD X55Y70VDD 25mOhm
L_X50Y70VDD_X60Y70VDD X55Y70VDD X60Y70VDD 2.91e-06nH
R_X50Y70VSS_X60Y70VSS X50Y70VSS X55Y70VSS 25mOhm
L_X50Y70VSS_X60Y70VSS X55Y70VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X70Y70VDD X60Y70VDD X65Y70VDD 25mOhm
L_X60Y70VDD_X70Y70VDD X65Y70VDD X70Y70VDD 2.91e-06nH
R_X60Y70VSS_X70Y70VSS X60Y70VSS X65Y70VSS 25mOhm
L_X60Y70VSS_X70Y70VSS X65Y70VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X80Y70VDD X70Y70VDD X75Y70VDD 25mOhm
L_X70Y70VDD_X80Y70VDD X75Y70VDD X80Y70VDD 2.91e-06nH
R_X70Y70VSS_X80Y70VSS X70Y70VSS X75Y70VSS 25mOhm
L_X70Y70VSS_X80Y70VSS X75Y70VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X90Y70VDD X80Y70VDD X85Y70VDD 25mOhm
L_X80Y70VDD_X90Y70VDD X85Y70VDD X90Y70VDD 2.91e-06nH
R_X80Y70VSS_X90Y70VSS X80Y70VSS X85Y70VSS 25mOhm
L_X80Y70VSS_X90Y70VSS X85Y70VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X100Y70VDD X90Y70VDD X95Y70VDD 25mOhm
L_X90Y70VDD_X100Y70VDD X95Y70VDD X100Y70VDD 2.91e-06nH
R_X90Y70VSS_X100Y70VSS X90Y70VSS X95Y70VSS 25mOhm
L_X90Y70VSS_X100Y70VSS X95Y70VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X110Y70VDD X100Y70VDD X105Y70VDD 25mOhm
L_X100Y70VDD_X110Y70VDD X105Y70VDD X110Y70VDD 2.91e-06nH
R_X100Y70VSS_X110Y70VSS X100Y70VSS X105Y70VSS 25mOhm
L_X100Y70VSS_X110Y70VSS X105Y70VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X120Y70VDD X110Y70VDD X115Y70VDD 25mOhm
L_X110Y70VDD_X120Y70VDD X115Y70VDD X120Y70VDD 2.91e-06nH
R_X110Y70VSS_X120Y70VSS X110Y70VSS X115Y70VSS 25mOhm
L_X110Y70VSS_X120Y70VSS X115Y70VSS X120Y70VSS 2.91e-06nH
R_X10Y80VDD_X20Y80VDD X10Y80VDD X15Y80VDD 25mOhm
L_X10Y80VDD_X20Y80VDD X15Y80VDD X20Y80VDD 2.91e-06nH
R_X10Y80VSS_X20Y80VSS X10Y80VSS X15Y80VSS 25mOhm
L_X10Y80VSS_X20Y80VSS X15Y80VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X30Y80VDD X20Y80VDD X25Y80VDD 25mOhm
L_X20Y80VDD_X30Y80VDD X25Y80VDD X30Y80VDD 2.91e-06nH
R_X20Y80VSS_X30Y80VSS X20Y80VSS X25Y80VSS 25mOhm
L_X20Y80VSS_X30Y80VSS X25Y80VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X40Y80VDD X30Y80VDD X35Y80VDD 25mOhm
L_X30Y80VDD_X40Y80VDD X35Y80VDD X40Y80VDD 2.91e-06nH
R_X30Y80VSS_X40Y80VSS X30Y80VSS X35Y80VSS 25mOhm
L_X30Y80VSS_X40Y80VSS X35Y80VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X50Y80VDD X40Y80VDD X45Y80VDD 25mOhm
L_X40Y80VDD_X50Y80VDD X45Y80VDD X50Y80VDD 2.91e-06nH
R_X40Y80VSS_X50Y80VSS X40Y80VSS X45Y80VSS 25mOhm
L_X40Y80VSS_X50Y80VSS X45Y80VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X60Y80VDD X50Y80VDD X55Y80VDD 25mOhm
L_X50Y80VDD_X60Y80VDD X55Y80VDD X60Y80VDD 2.91e-06nH
R_X50Y80VSS_X60Y80VSS X50Y80VSS X55Y80VSS 25mOhm
L_X50Y80VSS_X60Y80VSS X55Y80VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X70Y80VDD X60Y80VDD X65Y80VDD 25mOhm
L_X60Y80VDD_X70Y80VDD X65Y80VDD X70Y80VDD 2.91e-06nH
R_X60Y80VSS_X70Y80VSS X60Y80VSS X65Y80VSS 25mOhm
L_X60Y80VSS_X70Y80VSS X65Y80VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X80Y80VDD X70Y80VDD X75Y80VDD 25mOhm
L_X70Y80VDD_X80Y80VDD X75Y80VDD X80Y80VDD 2.91e-06nH
R_X70Y80VSS_X80Y80VSS X70Y80VSS X75Y80VSS 25mOhm
L_X70Y80VSS_X80Y80VSS X75Y80VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X90Y80VDD X80Y80VDD X85Y80VDD 25mOhm
L_X80Y80VDD_X90Y80VDD X85Y80VDD X90Y80VDD 2.91e-06nH
R_X80Y80VSS_X90Y80VSS X80Y80VSS X85Y80VSS 25mOhm
L_X80Y80VSS_X90Y80VSS X85Y80VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X100Y80VDD X90Y80VDD X95Y80VDD 25mOhm
L_X90Y80VDD_X100Y80VDD X95Y80VDD X100Y80VDD 2.91e-06nH
R_X90Y80VSS_X100Y80VSS X90Y80VSS X95Y80VSS 25mOhm
L_X90Y80VSS_X100Y80VSS X95Y80VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X110Y80VDD X100Y80VDD X105Y80VDD 25mOhm
L_X100Y80VDD_X110Y80VDD X105Y80VDD X110Y80VDD 2.91e-06nH
R_X100Y80VSS_X110Y80VSS X100Y80VSS X105Y80VSS 25mOhm
L_X100Y80VSS_X110Y80VSS X105Y80VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X120Y80VDD X110Y80VDD X115Y80VDD 25mOhm
L_X110Y80VDD_X120Y80VDD X115Y80VDD X120Y80VDD 2.91e-06nH
R_X110Y80VSS_X120Y80VSS X110Y80VSS X115Y80VSS 25mOhm
L_X110Y80VSS_X120Y80VSS X115Y80VSS X120Y80VSS 2.91e-06nH
R_X10Y90VDD_X20Y90VDD X10Y90VDD X15Y90VDD 25mOhm
L_X10Y90VDD_X20Y90VDD X15Y90VDD X20Y90VDD 2.91e-06nH
R_X10Y90VSS_X20Y90VSS X10Y90VSS X15Y90VSS 25mOhm
L_X10Y90VSS_X20Y90VSS X15Y90VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X30Y90VDD X20Y90VDD X25Y90VDD 25mOhm
L_X20Y90VDD_X30Y90VDD X25Y90VDD X30Y90VDD 2.91e-06nH
R_X20Y90VSS_X30Y90VSS X20Y90VSS X25Y90VSS 25mOhm
L_X20Y90VSS_X30Y90VSS X25Y90VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X40Y90VDD X30Y90VDD X35Y90VDD 25mOhm
L_X30Y90VDD_X40Y90VDD X35Y90VDD X40Y90VDD 2.91e-06nH
R_X30Y90VSS_X40Y90VSS X30Y90VSS X35Y90VSS 25mOhm
L_X30Y90VSS_X40Y90VSS X35Y90VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X50Y90VDD X40Y90VDD X45Y90VDD 25mOhm
L_X40Y90VDD_X50Y90VDD X45Y90VDD X50Y90VDD 2.91e-06nH
R_X40Y90VSS_X50Y90VSS X40Y90VSS X45Y90VSS 25mOhm
L_X40Y90VSS_X50Y90VSS X45Y90VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X60Y90VDD X50Y90VDD X55Y90VDD 25mOhm
L_X50Y90VDD_X60Y90VDD X55Y90VDD X60Y90VDD 2.91e-06nH
R_X50Y90VSS_X60Y90VSS X50Y90VSS X55Y90VSS 25mOhm
L_X50Y90VSS_X60Y90VSS X55Y90VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X70Y90VDD X60Y90VDD X65Y90VDD 25mOhm
L_X60Y90VDD_X70Y90VDD X65Y90VDD X70Y90VDD 2.91e-06nH
R_X60Y90VSS_X70Y90VSS X60Y90VSS X65Y90VSS 25mOhm
L_X60Y90VSS_X70Y90VSS X65Y90VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X80Y90VDD X70Y90VDD X75Y90VDD 25mOhm
L_X70Y90VDD_X80Y90VDD X75Y90VDD X80Y90VDD 2.91e-06nH
R_X70Y90VSS_X80Y90VSS X70Y90VSS X75Y90VSS 25mOhm
L_X70Y90VSS_X80Y90VSS X75Y90VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X90Y90VDD X80Y90VDD X85Y90VDD 25mOhm
L_X80Y90VDD_X90Y90VDD X85Y90VDD X90Y90VDD 2.91e-06nH
R_X80Y90VSS_X90Y90VSS X80Y90VSS X85Y90VSS 25mOhm
L_X80Y90VSS_X90Y90VSS X85Y90VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X100Y90VDD X90Y90VDD X95Y90VDD 25mOhm
L_X90Y90VDD_X100Y90VDD X95Y90VDD X100Y90VDD 2.91e-06nH
R_X90Y90VSS_X100Y90VSS X90Y90VSS X95Y90VSS 25mOhm
L_X90Y90VSS_X100Y90VSS X95Y90VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X110Y90VDD X100Y90VDD X105Y90VDD 25mOhm
L_X100Y90VDD_X110Y90VDD X105Y90VDD X110Y90VDD 2.91e-06nH
R_X100Y90VSS_X110Y90VSS X100Y90VSS X105Y90VSS 25mOhm
L_X100Y90VSS_X110Y90VSS X105Y90VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X120Y90VDD X110Y90VDD X115Y90VDD 25mOhm
L_X110Y90VDD_X120Y90VDD X115Y90VDD X120Y90VDD 2.91e-06nH
R_X110Y90VSS_X120Y90VSS X110Y90VSS X115Y90VSS 25mOhm
L_X110Y90VSS_X120Y90VSS X115Y90VSS X120Y90VSS 2.91e-06nH
R_X10Y100VDD_X20Y100VDD X10Y100VDD X15Y100VDD 25mOhm
L_X10Y100VDD_X20Y100VDD X15Y100VDD X20Y100VDD 2.91e-06nH
R_X10Y100VSS_X20Y100VSS X10Y100VSS X15Y100VSS 25mOhm
L_X10Y100VSS_X20Y100VSS X15Y100VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X30Y100VDD X20Y100VDD X25Y100VDD 25mOhm
L_X20Y100VDD_X30Y100VDD X25Y100VDD X30Y100VDD 2.91e-06nH
R_X20Y100VSS_X30Y100VSS X20Y100VSS X25Y100VSS 25mOhm
L_X20Y100VSS_X30Y100VSS X25Y100VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X40Y100VDD X30Y100VDD X35Y100VDD 25mOhm
L_X30Y100VDD_X40Y100VDD X35Y100VDD X40Y100VDD 2.91e-06nH
R_X30Y100VSS_X40Y100VSS X30Y100VSS X35Y100VSS 25mOhm
L_X30Y100VSS_X40Y100VSS X35Y100VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X50Y100VDD X40Y100VDD X45Y100VDD 25mOhm
L_X40Y100VDD_X50Y100VDD X45Y100VDD X50Y100VDD 2.91e-06nH
R_X40Y100VSS_X50Y100VSS X40Y100VSS X45Y100VSS 25mOhm
L_X40Y100VSS_X50Y100VSS X45Y100VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X60Y100VDD X50Y100VDD X55Y100VDD 25mOhm
L_X50Y100VDD_X60Y100VDD X55Y100VDD X60Y100VDD 2.91e-06nH
R_X50Y100VSS_X60Y100VSS X50Y100VSS X55Y100VSS 25mOhm
L_X50Y100VSS_X60Y100VSS X55Y100VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X70Y100VDD X60Y100VDD X65Y100VDD 25mOhm
L_X60Y100VDD_X70Y100VDD X65Y100VDD X70Y100VDD 2.91e-06nH
R_X60Y100VSS_X70Y100VSS X60Y100VSS X65Y100VSS 25mOhm
L_X60Y100VSS_X70Y100VSS X65Y100VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X80Y100VDD X70Y100VDD X75Y100VDD 25mOhm
L_X70Y100VDD_X80Y100VDD X75Y100VDD X80Y100VDD 2.91e-06nH
R_X70Y100VSS_X80Y100VSS X70Y100VSS X75Y100VSS 25mOhm
L_X70Y100VSS_X80Y100VSS X75Y100VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X90Y100VDD X80Y100VDD X85Y100VDD 25mOhm
L_X80Y100VDD_X90Y100VDD X85Y100VDD X90Y100VDD 2.91e-06nH
R_X80Y100VSS_X90Y100VSS X80Y100VSS X85Y100VSS 25mOhm
L_X80Y100VSS_X90Y100VSS X85Y100VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X100Y100VDD X90Y100VDD X95Y100VDD 25mOhm
L_X90Y100VDD_X100Y100VDD X95Y100VDD X100Y100VDD 2.91e-06nH
R_X90Y100VSS_X100Y100VSS X90Y100VSS X95Y100VSS 25mOhm
L_X90Y100VSS_X100Y100VSS X95Y100VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X110Y100VDD X100Y100VDD X105Y100VDD 25mOhm
L_X100Y100VDD_X110Y100VDD X105Y100VDD X110Y100VDD 2.91e-06nH
R_X100Y100VSS_X110Y100VSS X100Y100VSS X105Y100VSS 25mOhm
L_X100Y100VSS_X110Y100VSS X105Y100VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X120Y100VDD X110Y100VDD X115Y100VDD 25mOhm
L_X110Y100VDD_X120Y100VDD X115Y100VDD X120Y100VDD 2.91e-06nH
R_X110Y100VSS_X120Y100VSS X110Y100VSS X115Y100VSS 25mOhm
L_X110Y100VSS_X120Y100VSS X115Y100VSS X120Y100VSS 2.91e-06nH
R_X10Y110VDD_X20Y110VDD X10Y110VDD X15Y110VDD 25mOhm
L_X10Y110VDD_X20Y110VDD X15Y110VDD X20Y110VDD 2.91e-06nH
R_X10Y110VSS_X20Y110VSS X10Y110VSS X15Y110VSS 25mOhm
L_X10Y110VSS_X20Y110VSS X15Y110VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X30Y110VDD X20Y110VDD X25Y110VDD 25mOhm
L_X20Y110VDD_X30Y110VDD X25Y110VDD X30Y110VDD 2.91e-06nH
R_X20Y110VSS_X30Y110VSS X20Y110VSS X25Y110VSS 25mOhm
L_X20Y110VSS_X30Y110VSS X25Y110VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X40Y110VDD X30Y110VDD X35Y110VDD 25mOhm
L_X30Y110VDD_X40Y110VDD X35Y110VDD X40Y110VDD 2.91e-06nH
R_X30Y110VSS_X40Y110VSS X30Y110VSS X35Y110VSS 25mOhm
L_X30Y110VSS_X40Y110VSS X35Y110VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X50Y110VDD X40Y110VDD X45Y110VDD 25mOhm
L_X40Y110VDD_X50Y110VDD X45Y110VDD X50Y110VDD 2.91e-06nH
R_X40Y110VSS_X50Y110VSS X40Y110VSS X45Y110VSS 25mOhm
L_X40Y110VSS_X50Y110VSS X45Y110VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X60Y110VDD X50Y110VDD X55Y110VDD 25mOhm
L_X50Y110VDD_X60Y110VDD X55Y110VDD X60Y110VDD 2.91e-06nH
R_X50Y110VSS_X60Y110VSS X50Y110VSS X55Y110VSS 25mOhm
L_X50Y110VSS_X60Y110VSS X55Y110VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X70Y110VDD X60Y110VDD X65Y110VDD 25mOhm
L_X60Y110VDD_X70Y110VDD X65Y110VDD X70Y110VDD 2.91e-06nH
R_X60Y110VSS_X70Y110VSS X60Y110VSS X65Y110VSS 25mOhm
L_X60Y110VSS_X70Y110VSS X65Y110VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X80Y110VDD X70Y110VDD X75Y110VDD 25mOhm
L_X70Y110VDD_X80Y110VDD X75Y110VDD X80Y110VDD 2.91e-06nH
R_X70Y110VSS_X80Y110VSS X70Y110VSS X75Y110VSS 25mOhm
L_X70Y110VSS_X80Y110VSS X75Y110VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X90Y110VDD X80Y110VDD X85Y110VDD 25mOhm
L_X80Y110VDD_X90Y110VDD X85Y110VDD X90Y110VDD 2.91e-06nH
R_X80Y110VSS_X90Y110VSS X80Y110VSS X85Y110VSS 25mOhm
L_X80Y110VSS_X90Y110VSS X85Y110VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X100Y110VDD X90Y110VDD X95Y110VDD 25mOhm
L_X90Y110VDD_X100Y110VDD X95Y110VDD X100Y110VDD 2.91e-06nH
R_X90Y110VSS_X100Y110VSS X90Y110VSS X95Y110VSS 25mOhm
L_X90Y110VSS_X100Y110VSS X95Y110VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X110Y110VDD X100Y110VDD X105Y110VDD 25mOhm
L_X100Y110VDD_X110Y110VDD X105Y110VDD X110Y110VDD 2.91e-06nH
R_X100Y110VSS_X110Y110VSS X100Y110VSS X105Y110VSS 25mOhm
L_X100Y110VSS_X110Y110VSS X105Y110VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X120Y110VDD X110Y110VDD X115Y110VDD 25mOhm
L_X110Y110VDD_X120Y110VDD X115Y110VDD X120Y110VDD 2.91e-06nH
R_X110Y110VSS_X120Y110VSS X110Y110VSS X115Y110VSS 25mOhm
L_X110Y110VSS_X120Y110VSS X115Y110VSS X120Y110VSS 2.91e-06nH
R_X10Y120VDD_X20Y120VDD X10Y120VDD X15Y120VDD 25mOhm
L_X10Y120VDD_X20Y120VDD X15Y120VDD X20Y120VDD 2.91e-06nH
R_X10Y120VSS_X20Y120VSS X10Y120VSS X15Y120VSS 25mOhm
L_X10Y120VSS_X20Y120VSS X15Y120VSS X20Y120VSS 2.91e-06nH
R_X20Y120VDD_X30Y120VDD X20Y120VDD X25Y120VDD 25mOhm
L_X20Y120VDD_X30Y120VDD X25Y120VDD X30Y120VDD 2.91e-06nH
R_X20Y120VSS_X30Y120VSS X20Y120VSS X25Y120VSS 25mOhm
L_X20Y120VSS_X30Y120VSS X25Y120VSS X30Y120VSS 2.91e-06nH
R_X30Y120VDD_X40Y120VDD X30Y120VDD X35Y120VDD 25mOhm
L_X30Y120VDD_X40Y120VDD X35Y120VDD X40Y120VDD 2.91e-06nH
R_X30Y120VSS_X40Y120VSS X30Y120VSS X35Y120VSS 25mOhm
L_X30Y120VSS_X40Y120VSS X35Y120VSS X40Y120VSS 2.91e-06nH
R_X40Y120VDD_X50Y120VDD X40Y120VDD X45Y120VDD 25mOhm
L_X40Y120VDD_X50Y120VDD X45Y120VDD X50Y120VDD 2.91e-06nH
R_X40Y120VSS_X50Y120VSS X40Y120VSS X45Y120VSS 25mOhm
L_X40Y120VSS_X50Y120VSS X45Y120VSS X50Y120VSS 2.91e-06nH
R_X50Y120VDD_X60Y120VDD X50Y120VDD X55Y120VDD 25mOhm
L_X50Y120VDD_X60Y120VDD X55Y120VDD X60Y120VDD 2.91e-06nH
R_X50Y120VSS_X60Y120VSS X50Y120VSS X55Y120VSS 25mOhm
L_X50Y120VSS_X60Y120VSS X55Y120VSS X60Y120VSS 2.91e-06nH
R_X60Y120VDD_X70Y120VDD X60Y120VDD X65Y120VDD 25mOhm
L_X60Y120VDD_X70Y120VDD X65Y120VDD X70Y120VDD 2.91e-06nH
R_X60Y120VSS_X70Y120VSS X60Y120VSS X65Y120VSS 25mOhm
L_X60Y120VSS_X70Y120VSS X65Y120VSS X70Y120VSS 2.91e-06nH
R_X70Y120VDD_X80Y120VDD X70Y120VDD X75Y120VDD 25mOhm
L_X70Y120VDD_X80Y120VDD X75Y120VDD X80Y120VDD 2.91e-06nH
R_X70Y120VSS_X80Y120VSS X70Y120VSS X75Y120VSS 25mOhm
L_X70Y120VSS_X80Y120VSS X75Y120VSS X80Y120VSS 2.91e-06nH
R_X80Y120VDD_X90Y120VDD X80Y120VDD X85Y120VDD 25mOhm
L_X80Y120VDD_X90Y120VDD X85Y120VDD X90Y120VDD 2.91e-06nH
R_X80Y120VSS_X90Y120VSS X80Y120VSS X85Y120VSS 25mOhm
L_X80Y120VSS_X90Y120VSS X85Y120VSS X90Y120VSS 2.91e-06nH
R_X90Y120VDD_X100Y120VDD X90Y120VDD X95Y120VDD 25mOhm
L_X90Y120VDD_X100Y120VDD X95Y120VDD X100Y120VDD 2.91e-06nH
R_X90Y120VSS_X100Y120VSS X90Y120VSS X95Y120VSS 25mOhm
L_X90Y120VSS_X100Y120VSS X95Y120VSS X100Y120VSS 2.91e-06nH
R_X100Y120VDD_X110Y120VDD X100Y120VDD X105Y120VDD 25mOhm
L_X100Y120VDD_X110Y120VDD X105Y120VDD X110Y120VDD 2.91e-06nH
R_X100Y120VSS_X110Y120VSS X100Y120VSS X105Y120VSS 25mOhm
L_X100Y120VSS_X110Y120VSS X105Y120VSS X110Y120VSS 2.91e-06nH
R_X110Y120VDD_X120Y120VDD X110Y120VDD X115Y120VDD 25mOhm
L_X110Y120VDD_X120Y120VDD X115Y120VDD X120Y120VDD 2.91e-06nH
R_X110Y120VSS_X120Y120VSS X110Y120VSS X115Y120VSS 25mOhm
L_X110Y120VSS_X120Y120VSS X115Y120VSS X120Y120VSS 2.91e-06nH
R_X10Y10VDD_X10Y20VDD X10Y10VDD X10Y15VDD 25mOhm
L_X10Y10VDD_X10Y20VDD X10Y15VDD X10Y20VDD 2.91e-06nH
R_X10Y10VSS_X10Y20VSS X10Y10VSS X10Y15VSS 25mOhm
L_X10Y10VSS_X10Y20VSS X10Y15VSS X10Y20VSS 2.91e-06nH
R_X10Y20VDD_X10Y30VDD X10Y20VDD X10Y25VDD 25mOhm
L_X10Y20VDD_X10Y30VDD X10Y25VDD X10Y30VDD 2.91e-06nH
R_X10Y20VSS_X10Y30VSS X10Y20VSS X10Y25VSS 25mOhm
L_X10Y20VSS_X10Y30VSS X10Y25VSS X10Y30VSS 2.91e-06nH
R_X10Y30VDD_X10Y40VDD X10Y30VDD X10Y35VDD 25mOhm
L_X10Y30VDD_X10Y40VDD X10Y35VDD X10Y40VDD 2.91e-06nH
R_X10Y30VSS_X10Y40VSS X10Y30VSS X10Y35VSS 25mOhm
L_X10Y30VSS_X10Y40VSS X10Y35VSS X10Y40VSS 2.91e-06nH
R_X10Y40VDD_X10Y50VDD X10Y40VDD X10Y45VDD 25mOhm
L_X10Y40VDD_X10Y50VDD X10Y45VDD X10Y50VDD 2.91e-06nH
R_X10Y40VSS_X10Y50VSS X10Y40VSS X10Y45VSS 25mOhm
L_X10Y40VSS_X10Y50VSS X10Y45VSS X10Y50VSS 2.91e-06nH
R_X10Y50VDD_X10Y60VDD X10Y50VDD X10Y55VDD 25mOhm
L_X10Y50VDD_X10Y60VDD X10Y55VDD X10Y60VDD 2.91e-06nH
R_X10Y50VSS_X10Y60VSS X10Y50VSS X10Y55VSS 25mOhm
L_X10Y50VSS_X10Y60VSS X10Y55VSS X10Y60VSS 2.91e-06nH
R_X10Y60VDD_X10Y70VDD X10Y60VDD X10Y65VDD 25mOhm
L_X10Y60VDD_X10Y70VDD X10Y65VDD X10Y70VDD 2.91e-06nH
R_X10Y60VSS_X10Y70VSS X10Y60VSS X10Y65VSS 25mOhm
L_X10Y60VSS_X10Y70VSS X10Y65VSS X10Y70VSS 2.91e-06nH
R_X10Y70VDD_X10Y80VDD X10Y70VDD X10Y75VDD 25mOhm
L_X10Y70VDD_X10Y80VDD X10Y75VDD X10Y80VDD 2.91e-06nH
R_X10Y70VSS_X10Y80VSS X10Y70VSS X10Y75VSS 25mOhm
L_X10Y70VSS_X10Y80VSS X10Y75VSS X10Y80VSS 2.91e-06nH
R_X10Y80VDD_X10Y90VDD X10Y80VDD X10Y85VDD 25mOhm
L_X10Y80VDD_X10Y90VDD X10Y85VDD X10Y90VDD 2.91e-06nH
R_X10Y80VSS_X10Y90VSS X10Y80VSS X10Y85VSS 25mOhm
L_X10Y80VSS_X10Y90VSS X10Y85VSS X10Y90VSS 2.91e-06nH
R_X10Y90VDD_X10Y100VDD X10Y90VDD X10Y95VDD 25mOhm
L_X10Y90VDD_X10Y100VDD X10Y95VDD X10Y100VDD 2.91e-06nH
R_X10Y90VSS_X10Y100VSS X10Y90VSS X10Y95VSS 25mOhm
L_X10Y90VSS_X10Y100VSS X10Y95VSS X10Y100VSS 2.91e-06nH
R_X10Y100VDD_X10Y110VDD X10Y100VDD X10Y105VDD 25mOhm
L_X10Y100VDD_X10Y110VDD X10Y105VDD X10Y110VDD 2.91e-06nH
R_X10Y100VSS_X10Y110VSS X10Y100VSS X10Y105VSS 25mOhm
L_X10Y100VSS_X10Y110VSS X10Y105VSS X10Y110VSS 2.91e-06nH
R_X10Y110VDD_X10Y120VDD X10Y110VDD X10Y115VDD 25mOhm
L_X10Y110VDD_X10Y120VDD X10Y115VDD X10Y120VDD 2.91e-06nH
R_X10Y110VSS_X10Y120VSS X10Y110VSS X10Y115VSS 25mOhm
L_X10Y110VSS_X10Y120VSS X10Y115VSS X10Y120VSS 2.91e-06nH
R_X20Y10VDD_X20Y20VDD X20Y10VDD X20Y15VDD 25mOhm
L_X20Y10VDD_X20Y20VDD X20Y15VDD X20Y20VDD 2.91e-06nH
R_X20Y10VSS_X20Y20VSS X20Y10VSS X20Y15VSS 25mOhm
L_X20Y10VSS_X20Y20VSS X20Y15VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X20Y30VDD X20Y20VDD X20Y25VDD 25mOhm
L_X20Y20VDD_X20Y30VDD X20Y25VDD X20Y30VDD 2.91e-06nH
R_X20Y20VSS_X20Y30VSS X20Y20VSS X20Y25VSS 25mOhm
L_X20Y20VSS_X20Y30VSS X20Y25VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X20Y40VDD X20Y30VDD X20Y35VDD 25mOhm
L_X20Y30VDD_X20Y40VDD X20Y35VDD X20Y40VDD 2.91e-06nH
R_X20Y30VSS_X20Y40VSS X20Y30VSS X20Y35VSS 25mOhm
L_X20Y30VSS_X20Y40VSS X20Y35VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X20Y50VDD X20Y40VDD X20Y45VDD 25mOhm
L_X20Y40VDD_X20Y50VDD X20Y45VDD X20Y50VDD 2.91e-06nH
R_X20Y40VSS_X20Y50VSS X20Y40VSS X20Y45VSS 25mOhm
L_X20Y40VSS_X20Y50VSS X20Y45VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X20Y60VDD X20Y50VDD X20Y55VDD 25mOhm
L_X20Y50VDD_X20Y60VDD X20Y55VDD X20Y60VDD 2.91e-06nH
R_X20Y50VSS_X20Y60VSS X20Y50VSS X20Y55VSS 25mOhm
L_X20Y50VSS_X20Y60VSS X20Y55VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X20Y70VDD X20Y60VDD X20Y65VDD 25mOhm
L_X20Y60VDD_X20Y70VDD X20Y65VDD X20Y70VDD 2.91e-06nH
R_X20Y60VSS_X20Y70VSS X20Y60VSS X20Y65VSS 25mOhm
L_X20Y60VSS_X20Y70VSS X20Y65VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X20Y80VDD X20Y70VDD X20Y75VDD 25mOhm
L_X20Y70VDD_X20Y80VDD X20Y75VDD X20Y80VDD 2.91e-06nH
R_X20Y70VSS_X20Y80VSS X20Y70VSS X20Y75VSS 25mOhm
L_X20Y70VSS_X20Y80VSS X20Y75VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X20Y90VDD X20Y80VDD X20Y85VDD 25mOhm
L_X20Y80VDD_X20Y90VDD X20Y85VDD X20Y90VDD 2.91e-06nH
R_X20Y80VSS_X20Y90VSS X20Y80VSS X20Y85VSS 25mOhm
L_X20Y80VSS_X20Y90VSS X20Y85VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X20Y100VDD X20Y90VDD X20Y95VDD 25mOhm
L_X20Y90VDD_X20Y100VDD X20Y95VDD X20Y100VDD 2.91e-06nH
R_X20Y90VSS_X20Y100VSS X20Y90VSS X20Y95VSS 25mOhm
L_X20Y90VSS_X20Y100VSS X20Y95VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X20Y110VDD X20Y100VDD X20Y105VDD 25mOhm
L_X20Y100VDD_X20Y110VDD X20Y105VDD X20Y110VDD 2.91e-06nH
R_X20Y100VSS_X20Y110VSS X20Y100VSS X20Y105VSS 25mOhm
L_X20Y100VSS_X20Y110VSS X20Y105VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X20Y120VDD X20Y110VDD X20Y115VDD 25mOhm
L_X20Y110VDD_X20Y120VDD X20Y115VDD X20Y120VDD 2.91e-06nH
R_X20Y110VSS_X20Y120VSS X20Y110VSS X20Y115VSS 25mOhm
L_X20Y110VSS_X20Y120VSS X20Y115VSS X20Y120VSS 2.91e-06nH
R_X30Y10VDD_X30Y20VDD X30Y10VDD X30Y15VDD 25mOhm
L_X30Y10VDD_X30Y20VDD X30Y15VDD X30Y20VDD 2.91e-06nH
R_X30Y10VSS_X30Y20VSS X30Y10VSS X30Y15VSS 25mOhm
L_X30Y10VSS_X30Y20VSS X30Y15VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X30Y30VDD X30Y20VDD X30Y25VDD 25mOhm
L_X30Y20VDD_X30Y30VDD X30Y25VDD X30Y30VDD 2.91e-06nH
R_X30Y20VSS_X30Y30VSS X30Y20VSS X30Y25VSS 25mOhm
L_X30Y20VSS_X30Y30VSS X30Y25VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X30Y40VDD X30Y30VDD X30Y35VDD 25mOhm
L_X30Y30VDD_X30Y40VDD X30Y35VDD X30Y40VDD 2.91e-06nH
R_X30Y30VSS_X30Y40VSS X30Y30VSS X30Y35VSS 25mOhm
L_X30Y30VSS_X30Y40VSS X30Y35VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X30Y50VDD X30Y40VDD X30Y45VDD 25mOhm
L_X30Y40VDD_X30Y50VDD X30Y45VDD X30Y50VDD 2.91e-06nH
R_X30Y40VSS_X30Y50VSS X30Y40VSS X30Y45VSS 25mOhm
L_X30Y40VSS_X30Y50VSS X30Y45VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X30Y60VDD X30Y50VDD X30Y55VDD 25mOhm
L_X30Y50VDD_X30Y60VDD X30Y55VDD X30Y60VDD 2.91e-06nH
R_X30Y50VSS_X30Y60VSS X30Y50VSS X30Y55VSS 25mOhm
L_X30Y50VSS_X30Y60VSS X30Y55VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X30Y70VDD X30Y60VDD X30Y65VDD 25mOhm
L_X30Y60VDD_X30Y70VDD X30Y65VDD X30Y70VDD 2.91e-06nH
R_X30Y60VSS_X30Y70VSS X30Y60VSS X30Y65VSS 25mOhm
L_X30Y60VSS_X30Y70VSS X30Y65VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X30Y80VDD X30Y70VDD X30Y75VDD 25mOhm
L_X30Y70VDD_X30Y80VDD X30Y75VDD X30Y80VDD 2.91e-06nH
R_X30Y70VSS_X30Y80VSS X30Y70VSS X30Y75VSS 25mOhm
L_X30Y70VSS_X30Y80VSS X30Y75VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X30Y90VDD X30Y80VDD X30Y85VDD 25mOhm
L_X30Y80VDD_X30Y90VDD X30Y85VDD X30Y90VDD 2.91e-06nH
R_X30Y80VSS_X30Y90VSS X30Y80VSS X30Y85VSS 25mOhm
L_X30Y80VSS_X30Y90VSS X30Y85VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X30Y100VDD X30Y90VDD X30Y95VDD 25mOhm
L_X30Y90VDD_X30Y100VDD X30Y95VDD X30Y100VDD 2.91e-06nH
R_X30Y90VSS_X30Y100VSS X30Y90VSS X30Y95VSS 25mOhm
L_X30Y90VSS_X30Y100VSS X30Y95VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X30Y110VDD X30Y100VDD X30Y105VDD 25mOhm
L_X30Y100VDD_X30Y110VDD X30Y105VDD X30Y110VDD 2.91e-06nH
R_X30Y100VSS_X30Y110VSS X30Y100VSS X30Y105VSS 25mOhm
L_X30Y100VSS_X30Y110VSS X30Y105VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X30Y120VDD X30Y110VDD X30Y115VDD 25mOhm
L_X30Y110VDD_X30Y120VDD X30Y115VDD X30Y120VDD 2.91e-06nH
R_X30Y110VSS_X30Y120VSS X30Y110VSS X30Y115VSS 25mOhm
L_X30Y110VSS_X30Y120VSS X30Y115VSS X30Y120VSS 2.91e-06nH
R_X40Y10VDD_X40Y20VDD X40Y10VDD X40Y15VDD 25mOhm
L_X40Y10VDD_X40Y20VDD X40Y15VDD X40Y20VDD 2.91e-06nH
R_X40Y10VSS_X40Y20VSS X40Y10VSS X40Y15VSS 25mOhm
L_X40Y10VSS_X40Y20VSS X40Y15VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X40Y30VDD X40Y20VDD X40Y25VDD 25mOhm
L_X40Y20VDD_X40Y30VDD X40Y25VDD X40Y30VDD 2.91e-06nH
R_X40Y20VSS_X40Y30VSS X40Y20VSS X40Y25VSS 25mOhm
L_X40Y20VSS_X40Y30VSS X40Y25VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X40Y40VDD X40Y30VDD X40Y35VDD 25mOhm
L_X40Y30VDD_X40Y40VDD X40Y35VDD X40Y40VDD 2.91e-06nH
R_X40Y30VSS_X40Y40VSS X40Y30VSS X40Y35VSS 25mOhm
L_X40Y30VSS_X40Y40VSS X40Y35VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X40Y50VDD X40Y40VDD X40Y45VDD 25mOhm
L_X40Y40VDD_X40Y50VDD X40Y45VDD X40Y50VDD 2.91e-06nH
R_X40Y40VSS_X40Y50VSS X40Y40VSS X40Y45VSS 25mOhm
L_X40Y40VSS_X40Y50VSS X40Y45VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X40Y60VDD X40Y50VDD X40Y55VDD 25mOhm
L_X40Y50VDD_X40Y60VDD X40Y55VDD X40Y60VDD 2.91e-06nH
R_X40Y50VSS_X40Y60VSS X40Y50VSS X40Y55VSS 25mOhm
L_X40Y50VSS_X40Y60VSS X40Y55VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X40Y70VDD X40Y60VDD X40Y65VDD 25mOhm
L_X40Y60VDD_X40Y70VDD X40Y65VDD X40Y70VDD 2.91e-06nH
R_X40Y60VSS_X40Y70VSS X40Y60VSS X40Y65VSS 25mOhm
L_X40Y60VSS_X40Y70VSS X40Y65VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X40Y80VDD X40Y70VDD X40Y75VDD 25mOhm
L_X40Y70VDD_X40Y80VDD X40Y75VDD X40Y80VDD 2.91e-06nH
R_X40Y70VSS_X40Y80VSS X40Y70VSS X40Y75VSS 25mOhm
L_X40Y70VSS_X40Y80VSS X40Y75VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X40Y90VDD X40Y80VDD X40Y85VDD 25mOhm
L_X40Y80VDD_X40Y90VDD X40Y85VDD X40Y90VDD 2.91e-06nH
R_X40Y80VSS_X40Y90VSS X40Y80VSS X40Y85VSS 25mOhm
L_X40Y80VSS_X40Y90VSS X40Y85VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X40Y100VDD X40Y90VDD X40Y95VDD 25mOhm
L_X40Y90VDD_X40Y100VDD X40Y95VDD X40Y100VDD 2.91e-06nH
R_X40Y90VSS_X40Y100VSS X40Y90VSS X40Y95VSS 25mOhm
L_X40Y90VSS_X40Y100VSS X40Y95VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X40Y110VDD X40Y100VDD X40Y105VDD 25mOhm
L_X40Y100VDD_X40Y110VDD X40Y105VDD X40Y110VDD 2.91e-06nH
R_X40Y100VSS_X40Y110VSS X40Y100VSS X40Y105VSS 25mOhm
L_X40Y100VSS_X40Y110VSS X40Y105VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X40Y120VDD X40Y110VDD X40Y115VDD 25mOhm
L_X40Y110VDD_X40Y120VDD X40Y115VDD X40Y120VDD 2.91e-06nH
R_X40Y110VSS_X40Y120VSS X40Y110VSS X40Y115VSS 25mOhm
L_X40Y110VSS_X40Y120VSS X40Y115VSS X40Y120VSS 2.91e-06nH
R_X50Y10VDD_X50Y20VDD X50Y10VDD X50Y15VDD 25mOhm
L_X50Y10VDD_X50Y20VDD X50Y15VDD X50Y20VDD 2.91e-06nH
R_X50Y10VSS_X50Y20VSS X50Y10VSS X50Y15VSS 25mOhm
L_X50Y10VSS_X50Y20VSS X50Y15VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X50Y30VDD X50Y20VDD X50Y25VDD 25mOhm
L_X50Y20VDD_X50Y30VDD X50Y25VDD X50Y30VDD 2.91e-06nH
R_X50Y20VSS_X50Y30VSS X50Y20VSS X50Y25VSS 25mOhm
L_X50Y20VSS_X50Y30VSS X50Y25VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X50Y40VDD X50Y30VDD X50Y35VDD 25mOhm
L_X50Y30VDD_X50Y40VDD X50Y35VDD X50Y40VDD 2.91e-06nH
R_X50Y30VSS_X50Y40VSS X50Y30VSS X50Y35VSS 25mOhm
L_X50Y30VSS_X50Y40VSS X50Y35VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X50Y50VDD X50Y40VDD X50Y45VDD 25mOhm
L_X50Y40VDD_X50Y50VDD X50Y45VDD X50Y50VDD 2.91e-06nH
R_X50Y40VSS_X50Y50VSS X50Y40VSS X50Y45VSS 25mOhm
L_X50Y40VSS_X50Y50VSS X50Y45VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X50Y60VDD X50Y50VDD X50Y55VDD 25mOhm
L_X50Y50VDD_X50Y60VDD X50Y55VDD X50Y60VDD 2.91e-06nH
R_X50Y50VSS_X50Y60VSS X50Y50VSS X50Y55VSS 25mOhm
L_X50Y50VSS_X50Y60VSS X50Y55VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X50Y70VDD X50Y60VDD X50Y65VDD 25mOhm
L_X50Y60VDD_X50Y70VDD X50Y65VDD X50Y70VDD 2.91e-06nH
R_X50Y60VSS_X50Y70VSS X50Y60VSS X50Y65VSS 25mOhm
L_X50Y60VSS_X50Y70VSS X50Y65VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X50Y80VDD X50Y70VDD X50Y75VDD 25mOhm
L_X50Y70VDD_X50Y80VDD X50Y75VDD X50Y80VDD 2.91e-06nH
R_X50Y70VSS_X50Y80VSS X50Y70VSS X50Y75VSS 25mOhm
L_X50Y70VSS_X50Y80VSS X50Y75VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X50Y90VDD X50Y80VDD X50Y85VDD 25mOhm
L_X50Y80VDD_X50Y90VDD X50Y85VDD X50Y90VDD 2.91e-06nH
R_X50Y80VSS_X50Y90VSS X50Y80VSS X50Y85VSS 25mOhm
L_X50Y80VSS_X50Y90VSS X50Y85VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X50Y100VDD X50Y90VDD X50Y95VDD 25mOhm
L_X50Y90VDD_X50Y100VDD X50Y95VDD X50Y100VDD 2.91e-06nH
R_X50Y90VSS_X50Y100VSS X50Y90VSS X50Y95VSS 25mOhm
L_X50Y90VSS_X50Y100VSS X50Y95VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X50Y110VDD X50Y100VDD X50Y105VDD 25mOhm
L_X50Y100VDD_X50Y110VDD X50Y105VDD X50Y110VDD 2.91e-06nH
R_X50Y100VSS_X50Y110VSS X50Y100VSS X50Y105VSS 25mOhm
L_X50Y100VSS_X50Y110VSS X50Y105VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X50Y120VDD X50Y110VDD X50Y115VDD 25mOhm
L_X50Y110VDD_X50Y120VDD X50Y115VDD X50Y120VDD 2.91e-06nH
R_X50Y110VSS_X50Y120VSS X50Y110VSS X50Y115VSS 25mOhm
L_X50Y110VSS_X50Y120VSS X50Y115VSS X50Y120VSS 2.91e-06nH
R_X60Y10VDD_X60Y20VDD X60Y10VDD X60Y15VDD 25mOhm
L_X60Y10VDD_X60Y20VDD X60Y15VDD X60Y20VDD 2.91e-06nH
R_X60Y10VSS_X60Y20VSS X60Y10VSS X60Y15VSS 25mOhm
L_X60Y10VSS_X60Y20VSS X60Y15VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X60Y30VDD X60Y20VDD X60Y25VDD 25mOhm
L_X60Y20VDD_X60Y30VDD X60Y25VDD X60Y30VDD 2.91e-06nH
R_X60Y20VSS_X60Y30VSS X60Y20VSS X60Y25VSS 25mOhm
L_X60Y20VSS_X60Y30VSS X60Y25VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X60Y40VDD X60Y30VDD X60Y35VDD 25mOhm
L_X60Y30VDD_X60Y40VDD X60Y35VDD X60Y40VDD 2.91e-06nH
R_X60Y30VSS_X60Y40VSS X60Y30VSS X60Y35VSS 25mOhm
L_X60Y30VSS_X60Y40VSS X60Y35VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X60Y50VDD X60Y40VDD X60Y45VDD 25mOhm
L_X60Y40VDD_X60Y50VDD X60Y45VDD X60Y50VDD 2.91e-06nH
R_X60Y40VSS_X60Y50VSS X60Y40VSS X60Y45VSS 25mOhm
L_X60Y40VSS_X60Y50VSS X60Y45VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X60Y60VDD X60Y50VDD X60Y55VDD 25mOhm
L_X60Y50VDD_X60Y60VDD X60Y55VDD X60Y60VDD 2.91e-06nH
R_X60Y50VSS_X60Y60VSS X60Y50VSS X60Y55VSS 25mOhm
L_X60Y50VSS_X60Y60VSS X60Y55VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X60Y70VDD X60Y60VDD X60Y65VDD 25mOhm
L_X60Y60VDD_X60Y70VDD X60Y65VDD X60Y70VDD 2.91e-06nH
R_X60Y60VSS_X60Y70VSS X60Y60VSS X60Y65VSS 25mOhm
L_X60Y60VSS_X60Y70VSS X60Y65VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X60Y80VDD X60Y70VDD X60Y75VDD 25mOhm
L_X60Y70VDD_X60Y80VDD X60Y75VDD X60Y80VDD 2.91e-06nH
R_X60Y70VSS_X60Y80VSS X60Y70VSS X60Y75VSS 25mOhm
L_X60Y70VSS_X60Y80VSS X60Y75VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X60Y90VDD X60Y80VDD X60Y85VDD 25mOhm
L_X60Y80VDD_X60Y90VDD X60Y85VDD X60Y90VDD 2.91e-06nH
R_X60Y80VSS_X60Y90VSS X60Y80VSS X60Y85VSS 25mOhm
L_X60Y80VSS_X60Y90VSS X60Y85VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X60Y100VDD X60Y90VDD X60Y95VDD 25mOhm
L_X60Y90VDD_X60Y100VDD X60Y95VDD X60Y100VDD 2.91e-06nH
R_X60Y90VSS_X60Y100VSS X60Y90VSS X60Y95VSS 25mOhm
L_X60Y90VSS_X60Y100VSS X60Y95VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X60Y110VDD X60Y100VDD X60Y105VDD 25mOhm
L_X60Y100VDD_X60Y110VDD X60Y105VDD X60Y110VDD 2.91e-06nH
R_X60Y100VSS_X60Y110VSS X60Y100VSS X60Y105VSS 25mOhm
L_X60Y100VSS_X60Y110VSS X60Y105VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X60Y120VDD X60Y110VDD X60Y115VDD 25mOhm
L_X60Y110VDD_X60Y120VDD X60Y115VDD X60Y120VDD 2.91e-06nH
R_X60Y110VSS_X60Y120VSS X60Y110VSS X60Y115VSS 25mOhm
L_X60Y110VSS_X60Y120VSS X60Y115VSS X60Y120VSS 2.91e-06nH
R_X70Y10VDD_X70Y20VDD X70Y10VDD X70Y15VDD 25mOhm
L_X70Y10VDD_X70Y20VDD X70Y15VDD X70Y20VDD 2.91e-06nH
R_X70Y10VSS_X70Y20VSS X70Y10VSS X70Y15VSS 25mOhm
L_X70Y10VSS_X70Y20VSS X70Y15VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X70Y30VDD X70Y20VDD X70Y25VDD 25mOhm
L_X70Y20VDD_X70Y30VDD X70Y25VDD X70Y30VDD 2.91e-06nH
R_X70Y20VSS_X70Y30VSS X70Y20VSS X70Y25VSS 25mOhm
L_X70Y20VSS_X70Y30VSS X70Y25VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X70Y40VDD X70Y30VDD X70Y35VDD 25mOhm
L_X70Y30VDD_X70Y40VDD X70Y35VDD X70Y40VDD 2.91e-06nH
R_X70Y30VSS_X70Y40VSS X70Y30VSS X70Y35VSS 25mOhm
L_X70Y30VSS_X70Y40VSS X70Y35VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X70Y50VDD X70Y40VDD X70Y45VDD 25mOhm
L_X70Y40VDD_X70Y50VDD X70Y45VDD X70Y50VDD 2.91e-06nH
R_X70Y40VSS_X70Y50VSS X70Y40VSS X70Y45VSS 25mOhm
L_X70Y40VSS_X70Y50VSS X70Y45VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X70Y60VDD X70Y50VDD X70Y55VDD 25mOhm
L_X70Y50VDD_X70Y60VDD X70Y55VDD X70Y60VDD 2.91e-06nH
R_X70Y50VSS_X70Y60VSS X70Y50VSS X70Y55VSS 25mOhm
L_X70Y50VSS_X70Y60VSS X70Y55VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X70Y70VDD X70Y60VDD X70Y65VDD 25mOhm
L_X70Y60VDD_X70Y70VDD X70Y65VDD X70Y70VDD 2.91e-06nH
R_X70Y60VSS_X70Y70VSS X70Y60VSS X70Y65VSS 25mOhm
L_X70Y60VSS_X70Y70VSS X70Y65VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X70Y80VDD X70Y70VDD X70Y75VDD 25mOhm
L_X70Y70VDD_X70Y80VDD X70Y75VDD X70Y80VDD 2.91e-06nH
R_X70Y70VSS_X70Y80VSS X70Y70VSS X70Y75VSS 25mOhm
L_X70Y70VSS_X70Y80VSS X70Y75VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X70Y90VDD X70Y80VDD X70Y85VDD 25mOhm
L_X70Y80VDD_X70Y90VDD X70Y85VDD X70Y90VDD 2.91e-06nH
R_X70Y80VSS_X70Y90VSS X70Y80VSS X70Y85VSS 25mOhm
L_X70Y80VSS_X70Y90VSS X70Y85VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X70Y100VDD X70Y90VDD X70Y95VDD 25mOhm
L_X70Y90VDD_X70Y100VDD X70Y95VDD X70Y100VDD 2.91e-06nH
R_X70Y90VSS_X70Y100VSS X70Y90VSS X70Y95VSS 25mOhm
L_X70Y90VSS_X70Y100VSS X70Y95VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X70Y110VDD X70Y100VDD X70Y105VDD 25mOhm
L_X70Y100VDD_X70Y110VDD X70Y105VDD X70Y110VDD 2.91e-06nH
R_X70Y100VSS_X70Y110VSS X70Y100VSS X70Y105VSS 25mOhm
L_X70Y100VSS_X70Y110VSS X70Y105VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X70Y120VDD X70Y110VDD X70Y115VDD 25mOhm
L_X70Y110VDD_X70Y120VDD X70Y115VDD X70Y120VDD 2.91e-06nH
R_X70Y110VSS_X70Y120VSS X70Y110VSS X70Y115VSS 25mOhm
L_X70Y110VSS_X70Y120VSS X70Y115VSS X70Y120VSS 2.91e-06nH
R_X80Y10VDD_X80Y20VDD X80Y10VDD X80Y15VDD 25mOhm
L_X80Y10VDD_X80Y20VDD X80Y15VDD X80Y20VDD 2.91e-06nH
R_X80Y10VSS_X80Y20VSS X80Y10VSS X80Y15VSS 25mOhm
L_X80Y10VSS_X80Y20VSS X80Y15VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X80Y30VDD X80Y20VDD X80Y25VDD 25mOhm
L_X80Y20VDD_X80Y30VDD X80Y25VDD X80Y30VDD 2.91e-06nH
R_X80Y20VSS_X80Y30VSS X80Y20VSS X80Y25VSS 25mOhm
L_X80Y20VSS_X80Y30VSS X80Y25VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X80Y40VDD X80Y30VDD X80Y35VDD 25mOhm
L_X80Y30VDD_X80Y40VDD X80Y35VDD X80Y40VDD 2.91e-06nH
R_X80Y30VSS_X80Y40VSS X80Y30VSS X80Y35VSS 25mOhm
L_X80Y30VSS_X80Y40VSS X80Y35VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X80Y50VDD X80Y40VDD X80Y45VDD 25mOhm
L_X80Y40VDD_X80Y50VDD X80Y45VDD X80Y50VDD 2.91e-06nH
R_X80Y40VSS_X80Y50VSS X80Y40VSS X80Y45VSS 25mOhm
L_X80Y40VSS_X80Y50VSS X80Y45VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X80Y60VDD X80Y50VDD X80Y55VDD 25mOhm
L_X80Y50VDD_X80Y60VDD X80Y55VDD X80Y60VDD 2.91e-06nH
R_X80Y50VSS_X80Y60VSS X80Y50VSS X80Y55VSS 25mOhm
L_X80Y50VSS_X80Y60VSS X80Y55VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X80Y70VDD X80Y60VDD X80Y65VDD 25mOhm
L_X80Y60VDD_X80Y70VDD X80Y65VDD X80Y70VDD 2.91e-06nH
R_X80Y60VSS_X80Y70VSS X80Y60VSS X80Y65VSS 25mOhm
L_X80Y60VSS_X80Y70VSS X80Y65VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X80Y80VDD X80Y70VDD X80Y75VDD 25mOhm
L_X80Y70VDD_X80Y80VDD X80Y75VDD X80Y80VDD 2.91e-06nH
R_X80Y70VSS_X80Y80VSS X80Y70VSS X80Y75VSS 25mOhm
L_X80Y70VSS_X80Y80VSS X80Y75VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X80Y90VDD X80Y80VDD X80Y85VDD 25mOhm
L_X80Y80VDD_X80Y90VDD X80Y85VDD X80Y90VDD 2.91e-06nH
R_X80Y80VSS_X80Y90VSS X80Y80VSS X80Y85VSS 25mOhm
L_X80Y80VSS_X80Y90VSS X80Y85VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X80Y100VDD X80Y90VDD X80Y95VDD 25mOhm
L_X80Y90VDD_X80Y100VDD X80Y95VDD X80Y100VDD 2.91e-06nH
R_X80Y90VSS_X80Y100VSS X80Y90VSS X80Y95VSS 25mOhm
L_X80Y90VSS_X80Y100VSS X80Y95VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X80Y110VDD X80Y100VDD X80Y105VDD 25mOhm
L_X80Y100VDD_X80Y110VDD X80Y105VDD X80Y110VDD 2.91e-06nH
R_X80Y100VSS_X80Y110VSS X80Y100VSS X80Y105VSS 25mOhm
L_X80Y100VSS_X80Y110VSS X80Y105VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X80Y120VDD X80Y110VDD X80Y115VDD 25mOhm
L_X80Y110VDD_X80Y120VDD X80Y115VDD X80Y120VDD 2.91e-06nH
R_X80Y110VSS_X80Y120VSS X80Y110VSS X80Y115VSS 25mOhm
L_X80Y110VSS_X80Y120VSS X80Y115VSS X80Y120VSS 2.91e-06nH
R_X90Y10VDD_X90Y20VDD X90Y10VDD X90Y15VDD 25mOhm
L_X90Y10VDD_X90Y20VDD X90Y15VDD X90Y20VDD 2.91e-06nH
R_X90Y10VSS_X90Y20VSS X90Y10VSS X90Y15VSS 25mOhm
L_X90Y10VSS_X90Y20VSS X90Y15VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X90Y30VDD X90Y20VDD X90Y25VDD 25mOhm
L_X90Y20VDD_X90Y30VDD X90Y25VDD X90Y30VDD 2.91e-06nH
R_X90Y20VSS_X90Y30VSS X90Y20VSS X90Y25VSS 25mOhm
L_X90Y20VSS_X90Y30VSS X90Y25VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X90Y40VDD X90Y30VDD X90Y35VDD 25mOhm
L_X90Y30VDD_X90Y40VDD X90Y35VDD X90Y40VDD 2.91e-06nH
R_X90Y30VSS_X90Y40VSS X90Y30VSS X90Y35VSS 25mOhm
L_X90Y30VSS_X90Y40VSS X90Y35VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X90Y50VDD X90Y40VDD X90Y45VDD 25mOhm
L_X90Y40VDD_X90Y50VDD X90Y45VDD X90Y50VDD 2.91e-06nH
R_X90Y40VSS_X90Y50VSS X90Y40VSS X90Y45VSS 25mOhm
L_X90Y40VSS_X90Y50VSS X90Y45VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X90Y60VDD X90Y50VDD X90Y55VDD 25mOhm
L_X90Y50VDD_X90Y60VDD X90Y55VDD X90Y60VDD 2.91e-06nH
R_X90Y50VSS_X90Y60VSS X90Y50VSS X90Y55VSS 25mOhm
L_X90Y50VSS_X90Y60VSS X90Y55VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X90Y70VDD X90Y60VDD X90Y65VDD 25mOhm
L_X90Y60VDD_X90Y70VDD X90Y65VDD X90Y70VDD 2.91e-06nH
R_X90Y60VSS_X90Y70VSS X90Y60VSS X90Y65VSS 25mOhm
L_X90Y60VSS_X90Y70VSS X90Y65VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X90Y80VDD X90Y70VDD X90Y75VDD 25mOhm
L_X90Y70VDD_X90Y80VDD X90Y75VDD X90Y80VDD 2.91e-06nH
R_X90Y70VSS_X90Y80VSS X90Y70VSS X90Y75VSS 25mOhm
L_X90Y70VSS_X90Y80VSS X90Y75VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X90Y90VDD X90Y80VDD X90Y85VDD 25mOhm
L_X90Y80VDD_X90Y90VDD X90Y85VDD X90Y90VDD 2.91e-06nH
R_X90Y80VSS_X90Y90VSS X90Y80VSS X90Y85VSS 25mOhm
L_X90Y80VSS_X90Y90VSS X90Y85VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X90Y100VDD X90Y90VDD X90Y95VDD 25mOhm
L_X90Y90VDD_X90Y100VDD X90Y95VDD X90Y100VDD 2.91e-06nH
R_X90Y90VSS_X90Y100VSS X90Y90VSS X90Y95VSS 25mOhm
L_X90Y90VSS_X90Y100VSS X90Y95VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X90Y110VDD X90Y100VDD X90Y105VDD 25mOhm
L_X90Y100VDD_X90Y110VDD X90Y105VDD X90Y110VDD 2.91e-06nH
R_X90Y100VSS_X90Y110VSS X90Y100VSS X90Y105VSS 25mOhm
L_X90Y100VSS_X90Y110VSS X90Y105VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X90Y120VDD X90Y110VDD X90Y115VDD 25mOhm
L_X90Y110VDD_X90Y120VDD X90Y115VDD X90Y120VDD 2.91e-06nH
R_X90Y110VSS_X90Y120VSS X90Y110VSS X90Y115VSS 25mOhm
L_X90Y110VSS_X90Y120VSS X90Y115VSS X90Y120VSS 2.91e-06nH
R_X100Y10VDD_X100Y20VDD X100Y10VDD X100Y15VDD 25mOhm
L_X100Y10VDD_X100Y20VDD X100Y15VDD X100Y20VDD 2.91e-06nH
R_X100Y10VSS_X100Y20VSS X100Y10VSS X100Y15VSS 25mOhm
L_X100Y10VSS_X100Y20VSS X100Y15VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X100Y30VDD X100Y20VDD X100Y25VDD 25mOhm
L_X100Y20VDD_X100Y30VDD X100Y25VDD X100Y30VDD 2.91e-06nH
R_X100Y20VSS_X100Y30VSS X100Y20VSS X100Y25VSS 25mOhm
L_X100Y20VSS_X100Y30VSS X100Y25VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X100Y40VDD X100Y30VDD X100Y35VDD 25mOhm
L_X100Y30VDD_X100Y40VDD X100Y35VDD X100Y40VDD 2.91e-06nH
R_X100Y30VSS_X100Y40VSS X100Y30VSS X100Y35VSS 25mOhm
L_X100Y30VSS_X100Y40VSS X100Y35VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X100Y50VDD X100Y40VDD X100Y45VDD 25mOhm
L_X100Y40VDD_X100Y50VDD X100Y45VDD X100Y50VDD 2.91e-06nH
R_X100Y40VSS_X100Y50VSS X100Y40VSS X100Y45VSS 25mOhm
L_X100Y40VSS_X100Y50VSS X100Y45VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X100Y60VDD X100Y50VDD X100Y55VDD 25mOhm
L_X100Y50VDD_X100Y60VDD X100Y55VDD X100Y60VDD 2.91e-06nH
R_X100Y50VSS_X100Y60VSS X100Y50VSS X100Y55VSS 25mOhm
L_X100Y50VSS_X100Y60VSS X100Y55VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X100Y70VDD X100Y60VDD X100Y65VDD 25mOhm
L_X100Y60VDD_X100Y70VDD X100Y65VDD X100Y70VDD 2.91e-06nH
R_X100Y60VSS_X100Y70VSS X100Y60VSS X100Y65VSS 25mOhm
L_X100Y60VSS_X100Y70VSS X100Y65VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X100Y80VDD X100Y70VDD X100Y75VDD 25mOhm
L_X100Y70VDD_X100Y80VDD X100Y75VDD X100Y80VDD 2.91e-06nH
R_X100Y70VSS_X100Y80VSS X100Y70VSS X100Y75VSS 25mOhm
L_X100Y70VSS_X100Y80VSS X100Y75VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X100Y90VDD X100Y80VDD X100Y85VDD 25mOhm
L_X100Y80VDD_X100Y90VDD X100Y85VDD X100Y90VDD 2.91e-06nH
R_X100Y80VSS_X100Y90VSS X100Y80VSS X100Y85VSS 25mOhm
L_X100Y80VSS_X100Y90VSS X100Y85VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X100Y100VDD X100Y90VDD X100Y95VDD 25mOhm
L_X100Y90VDD_X100Y100VDD X100Y95VDD X100Y100VDD 2.91e-06nH
R_X100Y90VSS_X100Y100VSS X100Y90VSS X100Y95VSS 25mOhm
L_X100Y90VSS_X100Y100VSS X100Y95VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X100Y110VDD X100Y100VDD X100Y105VDD 25mOhm
L_X100Y100VDD_X100Y110VDD X100Y105VDD X100Y110VDD 2.91e-06nH
R_X100Y100VSS_X100Y110VSS X100Y100VSS X100Y105VSS 25mOhm
L_X100Y100VSS_X100Y110VSS X100Y105VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X100Y120VDD X100Y110VDD X100Y115VDD 25mOhm
L_X100Y110VDD_X100Y120VDD X100Y115VDD X100Y120VDD 2.91e-06nH
R_X100Y110VSS_X100Y120VSS X100Y110VSS X100Y115VSS 25mOhm
L_X100Y110VSS_X100Y120VSS X100Y115VSS X100Y120VSS 2.91e-06nH
R_X110Y10VDD_X110Y20VDD X110Y10VDD X110Y15VDD 25mOhm
L_X110Y10VDD_X110Y20VDD X110Y15VDD X110Y20VDD 2.91e-06nH
R_X110Y10VSS_X110Y20VSS X110Y10VSS X110Y15VSS 25mOhm
L_X110Y10VSS_X110Y20VSS X110Y15VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X110Y30VDD X110Y20VDD X110Y25VDD 25mOhm
L_X110Y20VDD_X110Y30VDD X110Y25VDD X110Y30VDD 2.91e-06nH
R_X110Y20VSS_X110Y30VSS X110Y20VSS X110Y25VSS 25mOhm
L_X110Y20VSS_X110Y30VSS X110Y25VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X110Y40VDD X110Y30VDD X110Y35VDD 25mOhm
L_X110Y30VDD_X110Y40VDD X110Y35VDD X110Y40VDD 2.91e-06nH
R_X110Y30VSS_X110Y40VSS X110Y30VSS X110Y35VSS 25mOhm
L_X110Y30VSS_X110Y40VSS X110Y35VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X110Y50VDD X110Y40VDD X110Y45VDD 25mOhm
L_X110Y40VDD_X110Y50VDD X110Y45VDD X110Y50VDD 2.91e-06nH
R_X110Y40VSS_X110Y50VSS X110Y40VSS X110Y45VSS 25mOhm
L_X110Y40VSS_X110Y50VSS X110Y45VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X110Y60VDD X110Y50VDD X110Y55VDD 25mOhm
L_X110Y50VDD_X110Y60VDD X110Y55VDD X110Y60VDD 2.91e-06nH
R_X110Y50VSS_X110Y60VSS X110Y50VSS X110Y55VSS 25mOhm
L_X110Y50VSS_X110Y60VSS X110Y55VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X110Y70VDD X110Y60VDD X110Y65VDD 25mOhm
L_X110Y60VDD_X110Y70VDD X110Y65VDD X110Y70VDD 2.91e-06nH
R_X110Y60VSS_X110Y70VSS X110Y60VSS X110Y65VSS 25mOhm
L_X110Y60VSS_X110Y70VSS X110Y65VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X110Y80VDD X110Y70VDD X110Y75VDD 25mOhm
L_X110Y70VDD_X110Y80VDD X110Y75VDD X110Y80VDD 2.91e-06nH
R_X110Y70VSS_X110Y80VSS X110Y70VSS X110Y75VSS 25mOhm
L_X110Y70VSS_X110Y80VSS X110Y75VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X110Y90VDD X110Y80VDD X110Y85VDD 25mOhm
L_X110Y80VDD_X110Y90VDD X110Y85VDD X110Y90VDD 2.91e-06nH
R_X110Y80VSS_X110Y90VSS X110Y80VSS X110Y85VSS 25mOhm
L_X110Y80VSS_X110Y90VSS X110Y85VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X110Y100VDD X110Y90VDD X110Y95VDD 25mOhm
L_X110Y90VDD_X110Y100VDD X110Y95VDD X110Y100VDD 2.91e-06nH
R_X110Y90VSS_X110Y100VSS X110Y90VSS X110Y95VSS 25mOhm
L_X110Y90VSS_X110Y100VSS X110Y95VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X110Y110VDD X110Y100VDD X110Y105VDD 25mOhm
L_X110Y100VDD_X110Y110VDD X110Y105VDD X110Y110VDD 2.91e-06nH
R_X110Y100VSS_X110Y110VSS X110Y100VSS X110Y105VSS 25mOhm
L_X110Y100VSS_X110Y110VSS X110Y105VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X110Y120VDD X110Y110VDD X110Y115VDD 25mOhm
L_X110Y110VDD_X110Y120VDD X110Y115VDD X110Y120VDD 2.91e-06nH
R_X110Y110VSS_X110Y120VSS X110Y110VSS X110Y115VSS 25mOhm
L_X110Y110VSS_X110Y120VSS X110Y115VSS X110Y120VSS 2.91e-06nH
R_X120Y10VDD_X120Y20VDD X120Y10VDD X120Y15VDD 25mOhm
L_X120Y10VDD_X120Y20VDD X120Y15VDD X120Y20VDD 2.91e-06nH
R_X120Y10VSS_X120Y20VSS X120Y10VSS X120Y15VSS 25mOhm
L_X120Y10VSS_X120Y20VSS X120Y15VSS X120Y20VSS 2.91e-06nH
R_X120Y20VDD_X120Y30VDD X120Y20VDD X120Y25VDD 25mOhm
L_X120Y20VDD_X120Y30VDD X120Y25VDD X120Y30VDD 2.91e-06nH
R_X120Y20VSS_X120Y30VSS X120Y20VSS X120Y25VSS 25mOhm
L_X120Y20VSS_X120Y30VSS X120Y25VSS X120Y30VSS 2.91e-06nH
R_X120Y30VDD_X120Y40VDD X120Y30VDD X120Y35VDD 25mOhm
L_X120Y30VDD_X120Y40VDD X120Y35VDD X120Y40VDD 2.91e-06nH
R_X120Y30VSS_X120Y40VSS X120Y30VSS X120Y35VSS 25mOhm
L_X120Y30VSS_X120Y40VSS X120Y35VSS X120Y40VSS 2.91e-06nH
R_X120Y40VDD_X120Y50VDD X120Y40VDD X120Y45VDD 25mOhm
L_X120Y40VDD_X120Y50VDD X120Y45VDD X120Y50VDD 2.91e-06nH
R_X120Y40VSS_X120Y50VSS X120Y40VSS X120Y45VSS 25mOhm
L_X120Y40VSS_X120Y50VSS X120Y45VSS X120Y50VSS 2.91e-06nH
R_X120Y50VDD_X120Y60VDD X120Y50VDD X120Y55VDD 25mOhm
L_X120Y50VDD_X120Y60VDD X120Y55VDD X120Y60VDD 2.91e-06nH
R_X120Y50VSS_X120Y60VSS X120Y50VSS X120Y55VSS 25mOhm
L_X120Y50VSS_X120Y60VSS X120Y55VSS X120Y60VSS 2.91e-06nH
R_X120Y60VDD_X120Y70VDD X120Y60VDD X120Y65VDD 25mOhm
L_X120Y60VDD_X120Y70VDD X120Y65VDD X120Y70VDD 2.91e-06nH
R_X120Y60VSS_X120Y70VSS X120Y60VSS X120Y65VSS 25mOhm
L_X120Y60VSS_X120Y70VSS X120Y65VSS X120Y70VSS 2.91e-06nH
R_X120Y70VDD_X120Y80VDD X120Y70VDD X120Y75VDD 25mOhm
L_X120Y70VDD_X120Y80VDD X120Y75VDD X120Y80VDD 2.91e-06nH
R_X120Y70VSS_X120Y80VSS X120Y70VSS X120Y75VSS 25mOhm
L_X120Y70VSS_X120Y80VSS X120Y75VSS X120Y80VSS 2.91e-06nH
R_X120Y80VDD_X120Y90VDD X120Y80VDD X120Y85VDD 25mOhm
L_X120Y80VDD_X120Y90VDD X120Y85VDD X120Y90VDD 2.91e-06nH
R_X120Y80VSS_X120Y90VSS X120Y80VSS X120Y85VSS 25mOhm
L_X120Y80VSS_X120Y90VSS X120Y85VSS X120Y90VSS 2.91e-06nH
R_X120Y90VDD_X120Y100VDD X120Y90VDD X120Y95VDD 25mOhm
L_X120Y90VDD_X120Y100VDD X120Y95VDD X120Y100VDD 2.91e-06nH
R_X120Y90VSS_X120Y100VSS X120Y90VSS X120Y95VSS 25mOhm
L_X120Y90VSS_X120Y100VSS X120Y95VSS X120Y100VSS 2.91e-06nH
R_X120Y100VDD_X120Y110VDD X120Y100VDD X120Y105VDD 25mOhm
L_X120Y100VDD_X120Y110VDD X120Y105VDD X120Y110VDD 2.91e-06nH
R_X120Y100VSS_X120Y110VSS X120Y100VSS X120Y105VSS 25mOhm
L_X120Y100VSS_X120Y110VSS X120Y105VSS X120Y110VSS 2.91e-06nH
R_X120Y110VDD_X120Y120VDD X120Y110VDD X120Y115VDD 25mOhm
L_X120Y110VDD_X120Y120VDD X120Y115VDD X120Y120VDD 2.91e-06nH
R_X120Y110VSS_X120Y120VSS X120Y110VSS X120Y115VSS 25mOhm
L_X120Y110VSS_X120Y120VSS X120Y115VSS X120Y120VSS 2.91e-06nH
C_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VSS 10nF
C_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VSS 10nF
C_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VSS 10nF
C_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VSS 10nF
C_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VSS 10nF
C_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VSS 10nF
C_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VSS 10nF
C_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VSS 10nF
C_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VSS 10nF
C_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VSS 10nF
C_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VSS 10nF
C_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VSS 10nF
C_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VSS 10nF
C_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VSS 10nF
C_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VSS 10nF
C_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VSS 10nF
C_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VSS 10nF
C_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VSS 10nF
C_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VSS 10nF
C_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VSS 10nF
C_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VSS 10nF
C_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VSS 10nF
C_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VSS 10nF
C_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VSS 10nF
C_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VSS 10nF
C_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VSS 10nF
C_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VSS 10nF
C_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VSS 10nF
C_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VSS 10nF
C_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VSS 10nF
C_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VSS 10nF
C_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VSS 10nF
C_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VSS 10nF
C_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VSS 10nF
C_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VSS 10nF
C_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VSS 10nF
C_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VSS 10nF
C_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VSS 10nF
C_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VSS 10nF
C_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VSS 10nF
C_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VSS 10nF
C_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VSS 10nF
C_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VSS 10nF
C_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VSS 10nF
C_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VSS 10nF
C_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VSS 10nF
C_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VSS 10nF
C_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VSS 10nF
C_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VSS 10nF
C_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VSS 10nF
C_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VSS 10nF
C_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VSS 10nF
C_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VSS 10nF
C_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VSS 10nF
C_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VSS 10nF
C_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VSS 10nF
C_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VSS 10nF
C_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VSS 10nF
C_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VSS 10nF
C_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VSS 10nF
C_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VSS 10nF
C_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VSS 10nF
C_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VSS 10nF
C_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VSS 10nF
C_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VSS 10nF
C_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VSS 10nF
C_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VSS 10nF
C_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VSS 10nF
C_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VSS 10nF
C_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VSS 10nF
C_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VSS 10nF
C_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VSS 10nF
C_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VSS 10nF
C_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VSS 10nF
C_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VSS 10nF
C_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VSS 10nF
C_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VSS 10nF
C_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VSS 10nF
C_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VSS 10nF
C_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VSS 10nF
C_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VSS 10nF
C_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VSS 10nF
C_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VSS 10nF
C_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VSS 10nF
C_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VSS 10nF
C_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VSS 10nF
C_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VSS 10nF
C_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VSS 10nF
C_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VSS 10nF
C_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VSS 10nF
C_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VSS 10nF
C_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VSS 10nF
C_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VSS 10nF
C_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VSS 10nF
C_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VSS 10nF
C_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VSS 10nF
C_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VSS 10nF
C_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VSS 10nF
C_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VSS 10nF
C_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VSS 10nF
C_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VSS 10nF
C_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VSS 10nF
C_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VSS 10nF
C_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VSS 10nF
C_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VSS 10nF
C_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VSS 10nF
C_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VSS 10nF
C_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VSS 10nF
C_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VSS 10nF
C_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VSS 10nF
C_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VSS 10nF
C_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VSS 10nF
C_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VSS 10nF
C_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VSS 10nF
C_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VSS 10nF
C_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VSS 10nF
C_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VSS 10nF
C_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VSS 10nF
C_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VSS 10nF
C_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VSS 10nF
C_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VSS 10nF
C_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VSS 10nF
C_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VSS 10nF
C_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VSS 10nF
C_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VSS 10nF
C_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VSS 10nF
C_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VSS 10nF
C_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VSS 10nF
C_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VSS 10nF
C_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VSS 10nF
C_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VSS 10nF
C_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VSS 10nF
C_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VSS 10nF
C_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VSS 10nF
C_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VSS 10nF
C_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VSS 10nF
C_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VSS 10nF
C_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VSS 10nF
C_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VSS 10nF
C_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VSS 10nF
C_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VSS 10nF
C_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VSS 10nF
C_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VSS 10nF
C_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VSS 10nF
I_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VDDDM 0.8 AC=1
V_X120Y120VDD_X120Y120VSS X120Y120VDDDM X120Y120VSS 0
I_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VDDDM 0.8 AC=1
V_X120Y10VDD_X120Y10VSS X120Y10VDDDM X120Y10VSS 0
I_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VDDDM 0.8 AC=1
V_X120Y20VDD_X120Y20VSS X120Y20VDDDM X120Y20VSS 0
I_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VDDDM 0.8 AC=1
V_X120Y30VDD_X120Y30VSS X120Y30VDDDM X120Y30VSS 0
I_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VDDDM 0.8 AC=1
V_X120Y40VDD_X120Y40VSS X120Y40VDDDM X120Y40VSS 0
I_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VDDDM 0.8 AC=1
V_X120Y50VDD_X120Y50VSS X120Y50VDDDM X120Y50VSS 0
I_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VDDDM 0.8 AC=1
V_X120Y60VDD_X120Y60VSS X120Y60VDDDM X120Y60VSS 0
I_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VDDDM 0.8 AC=1
V_X120Y70VDD_X120Y70VSS X120Y70VDDDM X120Y70VSS 0
I_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VDDDM 0.8 AC=1
V_X120Y80VDD_X120Y80VSS X120Y80VDDDM X120Y80VSS 0
I_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VDDDM 0.8 AC=1
V_X120Y90VDD_X120Y90VSS X120Y90VDDDM X120Y90VSS 0
I_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VDDDM 0.8 AC=1
V_X120Y100VDD_X120Y100VSS X120Y100VDDDM X120Y100VSS 0
I_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VDDDM 0.8 AC=1
V_X120Y110VDD_X120Y110VSS X120Y110VDDDM X120Y110VSS 0
I_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VDDDM 0.8 AC=1
V_X10Y120VDD_X10Y120VSS X10Y120VDDDM X10Y120VSS 0
I_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VDDDM 0.8 AC=1
V_X10Y10VDD_X10Y10VSS X10Y10VDDDM X10Y10VSS 0
I_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VDDDM 0.8 AC=1
V_X10Y20VDD_X10Y20VSS X10Y20VDDDM X10Y20VSS 0
I_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VDDDM 0.8 AC=1
V_X10Y30VDD_X10Y30VSS X10Y30VDDDM X10Y30VSS 0
I_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VDDDM 0.8 AC=1
V_X10Y40VDD_X10Y40VSS X10Y40VDDDM X10Y40VSS 0
I_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VDDDM 0.8 AC=1
V_X10Y50VDD_X10Y50VSS X10Y50VDDDM X10Y50VSS 0
I_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VDDDM 0.8 AC=1
V_X10Y60VDD_X10Y60VSS X10Y60VDDDM X10Y60VSS 0
I_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VDDDM 0.8 AC=1
V_X10Y70VDD_X10Y70VSS X10Y70VDDDM X10Y70VSS 0
I_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VDDDM 0.8 AC=1
V_X10Y80VDD_X10Y80VSS X10Y80VDDDM X10Y80VSS 0
I_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VDDDM 0.8 AC=1
V_X10Y90VDD_X10Y90VSS X10Y90VDDDM X10Y90VSS 0
I_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VDDDM 0.8 AC=1
V_X10Y100VDD_X10Y100VSS X10Y100VDDDM X10Y100VSS 0
I_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VDDDM 0.8 AC=1
V_X10Y110VDD_X10Y110VSS X10Y110VDDDM X10Y110VSS 0
I_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VDDDM 0.8 AC=1
V_X20Y120VDD_X20Y120VSS X20Y120VDDDM X20Y120VSS 0
I_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VDDDM 0.8 AC=1
V_X20Y10VDD_X20Y10VSS X20Y10VDDDM X20Y10VSS 0
I_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VDDDM 0.8 AC=1
V_X20Y20VDD_X20Y20VSS X20Y20VDDDM X20Y20VSS 0
I_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VDDDM 0.8 AC=1
V_X20Y30VDD_X20Y30VSS X20Y30VDDDM X20Y30VSS 0
I_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VDDDM 0.8 AC=1
V_X20Y40VDD_X20Y40VSS X20Y40VDDDM X20Y40VSS 0
I_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VDDDM 0.8 AC=1
V_X20Y50VDD_X20Y50VSS X20Y50VDDDM X20Y50VSS 0
I_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VDDDM 0.8 AC=1
V_X20Y60VDD_X20Y60VSS X20Y60VDDDM X20Y60VSS 0
I_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VDDDM 0.8 AC=1
V_X20Y70VDD_X20Y70VSS X20Y70VDDDM X20Y70VSS 0
I_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VDDDM 0.8 AC=1
V_X20Y80VDD_X20Y80VSS X20Y80VDDDM X20Y80VSS 0
I_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VDDDM 0.8 AC=1
V_X20Y90VDD_X20Y90VSS X20Y90VDDDM X20Y90VSS 0
I_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VDDDM 0.8 AC=1
V_X20Y100VDD_X20Y100VSS X20Y100VDDDM X20Y100VSS 0
I_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VDDDM 0.8 AC=1
V_X20Y110VDD_X20Y110VSS X20Y110VDDDM X20Y110VSS 0
I_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VDDDM 0.8 AC=1
V_X30Y120VDD_X30Y120VSS X30Y120VDDDM X30Y120VSS 0
I_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VDDDM 0.8 AC=1
V_X30Y10VDD_X30Y10VSS X30Y10VDDDM X30Y10VSS 0
I_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VDDDM 0.8 AC=1
V_X30Y20VDD_X30Y20VSS X30Y20VDDDM X30Y20VSS 0
I_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VDDDM 0.8 AC=1
V_X30Y30VDD_X30Y30VSS X30Y30VDDDM X30Y30VSS 0
I_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VDDDM 0.8 AC=1
V_X30Y40VDD_X30Y40VSS X30Y40VDDDM X30Y40VSS 0
I_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VDDDM 0.8 AC=1
V_X30Y50VDD_X30Y50VSS X30Y50VDDDM X30Y50VSS 0
I_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VDDDM 0.8 AC=1
V_X30Y60VDD_X30Y60VSS X30Y60VDDDM X30Y60VSS 0
I_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VDDDM 0.8 AC=1
V_X30Y70VDD_X30Y70VSS X30Y70VDDDM X30Y70VSS 0
I_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VDDDM 0.8 AC=1
V_X30Y80VDD_X30Y80VSS X30Y80VDDDM X30Y80VSS 0
I_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VDDDM 0.8 AC=1
V_X30Y90VDD_X30Y90VSS X30Y90VDDDM X30Y90VSS 0
I_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VDDDM 0.8 AC=1
V_X30Y100VDD_X30Y100VSS X30Y100VDDDM X30Y100VSS 0
I_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VDDDM 0.8 AC=1
V_X30Y110VDD_X30Y110VSS X30Y110VDDDM X30Y110VSS 0
I_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VDDDM 0.8 AC=1
V_X40Y120VDD_X40Y120VSS X40Y120VDDDM X40Y120VSS 0
I_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VDDDM 0.8 AC=1
V_X40Y10VDD_X40Y10VSS X40Y10VDDDM X40Y10VSS 0
I_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VDDDM 0.8 AC=1
V_X40Y20VDD_X40Y20VSS X40Y20VDDDM X40Y20VSS 0
I_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VDDDM 0.8 AC=1
V_X40Y30VDD_X40Y30VSS X40Y30VDDDM X40Y30VSS 0
I_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VDDDM 0.8 AC=1
V_X40Y40VDD_X40Y40VSS X40Y40VDDDM X40Y40VSS 0
I_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VDDDM 0.8 AC=1
V_X40Y50VDD_X40Y50VSS X40Y50VDDDM X40Y50VSS 0
I_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VDDDM 0.8 AC=1
V_X40Y60VDD_X40Y60VSS X40Y60VDDDM X40Y60VSS 0
I_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VDDDM 0.8 AC=1
V_X40Y70VDD_X40Y70VSS X40Y70VDDDM X40Y70VSS 0
I_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VDDDM 0.8 AC=1
V_X40Y80VDD_X40Y80VSS X40Y80VDDDM X40Y80VSS 0
I_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VDDDM 0.8 AC=1
V_X40Y90VDD_X40Y90VSS X40Y90VDDDM X40Y90VSS 0
I_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VDDDM 0.8 AC=1
V_X40Y100VDD_X40Y100VSS X40Y100VDDDM X40Y100VSS 0
I_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VDDDM 0.8 AC=1
V_X40Y110VDD_X40Y110VSS X40Y110VDDDM X40Y110VSS 0
I_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VDDDM 0.8 AC=1
V_X50Y120VDD_X50Y120VSS X50Y120VDDDM X50Y120VSS 0
I_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VDDDM 0.8 AC=1
V_X50Y10VDD_X50Y10VSS X50Y10VDDDM X50Y10VSS 0
I_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VDDDM 0.8 AC=1
V_X50Y20VDD_X50Y20VSS X50Y20VDDDM X50Y20VSS 0
I_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VDDDM 0.8 AC=1
V_X50Y30VDD_X50Y30VSS X50Y30VDDDM X50Y30VSS 0
I_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VDDDM 0.8 AC=1
V_X50Y40VDD_X50Y40VSS X50Y40VDDDM X50Y40VSS 0
I_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VDDDM 0.8 AC=1
V_X50Y50VDD_X50Y50VSS X50Y50VDDDM X50Y50VSS 0
I_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VDDDM 0.8 AC=1
V_X50Y60VDD_X50Y60VSS X50Y60VDDDM X50Y60VSS 0
I_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VDDDM 0.8 AC=1
V_X50Y70VDD_X50Y70VSS X50Y70VDDDM X50Y70VSS 0
I_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VDDDM 0.8 AC=1
V_X50Y80VDD_X50Y80VSS X50Y80VDDDM X50Y80VSS 0
I_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VDDDM 0.8 AC=1
V_X50Y90VDD_X50Y90VSS X50Y90VDDDM X50Y90VSS 0
I_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VDDDM 0.8 AC=1
V_X50Y100VDD_X50Y100VSS X50Y100VDDDM X50Y100VSS 0
I_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VDDDM 0.8 AC=1
V_X50Y110VDD_X50Y110VSS X50Y110VDDDM X50Y110VSS 0
I_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VDDDM 0.8 AC=1
V_X60Y120VDD_X60Y120VSS X60Y120VDDDM X60Y120VSS 0
I_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VDDDM 0.8 AC=1
V_X60Y10VDD_X60Y10VSS X60Y10VDDDM X60Y10VSS 0
I_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VDDDM 0.8 AC=1
V_X60Y20VDD_X60Y20VSS X60Y20VDDDM X60Y20VSS 0
I_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VDDDM 0.8 AC=1
V_X60Y30VDD_X60Y30VSS X60Y30VDDDM X60Y30VSS 0
I_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VDDDM 0.8 AC=1
V_X60Y40VDD_X60Y40VSS X60Y40VDDDM X60Y40VSS 0
I_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VDDDM 0.8 AC=1
V_X60Y50VDD_X60Y50VSS X60Y50VDDDM X60Y50VSS 0
I_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VDDDM 0.8 AC=1
V_X60Y60VDD_X60Y60VSS X60Y60VDDDM X60Y60VSS 0
I_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VDDDM 0.8 AC=1
V_X60Y70VDD_X60Y70VSS X60Y70VDDDM X60Y70VSS 0
I_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VDDDM 0.8 AC=1
V_X60Y80VDD_X60Y80VSS X60Y80VDDDM X60Y80VSS 0
I_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VDDDM 0.8 AC=1
V_X60Y90VDD_X60Y90VSS X60Y90VDDDM X60Y90VSS 0
I_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VDDDM 0.8 AC=1
V_X60Y100VDD_X60Y100VSS X60Y100VDDDM X60Y100VSS 0
I_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VDDDM 0.8 AC=1
V_X60Y110VDD_X60Y110VSS X60Y110VDDDM X60Y110VSS 0
I_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VDDDM 0.8 AC=1
V_X70Y120VDD_X70Y120VSS X70Y120VDDDM X70Y120VSS 0
I_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VDDDM 0.8 AC=1
V_X70Y10VDD_X70Y10VSS X70Y10VDDDM X70Y10VSS 0
I_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VDDDM 0.8 AC=1
V_X70Y20VDD_X70Y20VSS X70Y20VDDDM X70Y20VSS 0
I_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VDDDM 0.8 AC=1
V_X70Y30VDD_X70Y30VSS X70Y30VDDDM X70Y30VSS 0
I_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VDDDM 0.8 AC=1
V_X70Y40VDD_X70Y40VSS X70Y40VDDDM X70Y40VSS 0
I_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VDDDM 0.8 AC=1
V_X70Y50VDD_X70Y50VSS X70Y50VDDDM X70Y50VSS 0
I_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VDDDM 0.8 AC=1
V_X70Y60VDD_X70Y60VSS X70Y60VDDDM X70Y60VSS 0
I_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VDDDM 0.8 AC=1
V_X70Y70VDD_X70Y70VSS X70Y70VDDDM X70Y70VSS 0
I_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VDDDM 0.8 AC=1
V_X70Y80VDD_X70Y80VSS X70Y80VDDDM X70Y80VSS 0
I_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VDDDM 0.8 AC=1
V_X70Y90VDD_X70Y90VSS X70Y90VDDDM X70Y90VSS 0
I_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VDDDM 0.8 AC=1
V_X70Y100VDD_X70Y100VSS X70Y100VDDDM X70Y100VSS 0
I_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VDDDM 0.8 AC=1
V_X70Y110VDD_X70Y110VSS X70Y110VDDDM X70Y110VSS 0
I_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VDDDM 0.8 AC=1
V_X80Y120VDD_X80Y120VSS X80Y120VDDDM X80Y120VSS 0
I_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VDDDM 0.8 AC=1
V_X80Y10VDD_X80Y10VSS X80Y10VDDDM X80Y10VSS 0
I_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VDDDM 0.8 AC=1
V_X80Y20VDD_X80Y20VSS X80Y20VDDDM X80Y20VSS 0
I_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VDDDM 0.8 AC=1
V_X80Y30VDD_X80Y30VSS X80Y30VDDDM X80Y30VSS 0
I_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VDDDM 0.8 AC=1
V_X80Y40VDD_X80Y40VSS X80Y40VDDDM X80Y40VSS 0
I_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VDDDM 0.8 AC=1
V_X80Y50VDD_X80Y50VSS X80Y50VDDDM X80Y50VSS 0
I_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VDDDM 0.8 AC=1
V_X80Y60VDD_X80Y60VSS X80Y60VDDDM X80Y60VSS 0
I_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VDDDM 0.8 AC=1
V_X80Y70VDD_X80Y70VSS X80Y70VDDDM X80Y70VSS 0
I_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VDDDM 0.8 AC=1
V_X80Y80VDD_X80Y80VSS X80Y80VDDDM X80Y80VSS 0
I_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VDDDM 0.8 AC=1
V_X80Y90VDD_X80Y90VSS X80Y90VDDDM X80Y90VSS 0
I_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VDDDM 0.8 AC=1
V_X80Y100VDD_X80Y100VSS X80Y100VDDDM X80Y100VSS 0
I_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VDDDM 0.8 AC=1
V_X80Y110VDD_X80Y110VSS X80Y110VDDDM X80Y110VSS 0
I_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VDDDM 0.8 AC=1
V_X90Y120VDD_X90Y120VSS X90Y120VDDDM X90Y120VSS 0
I_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VDDDM 0.8 AC=1
V_X90Y10VDD_X90Y10VSS X90Y10VDDDM X90Y10VSS 0
I_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VDDDM 0.8 AC=1
V_X90Y20VDD_X90Y20VSS X90Y20VDDDM X90Y20VSS 0
I_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VDDDM 0.8 AC=1
V_X90Y30VDD_X90Y30VSS X90Y30VDDDM X90Y30VSS 0
I_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VDDDM 0.8 AC=1
V_X90Y40VDD_X90Y40VSS X90Y40VDDDM X90Y40VSS 0
I_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VDDDM 0.8 AC=1
V_X90Y50VDD_X90Y50VSS X90Y50VDDDM X90Y50VSS 0
I_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VDDDM 0.8 AC=1
V_X90Y60VDD_X90Y60VSS X90Y60VDDDM X90Y60VSS 0
I_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VDDDM 0.8 AC=1
V_X90Y70VDD_X90Y70VSS X90Y70VDDDM X90Y70VSS 0
I_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VDDDM 0.8 AC=1
V_X90Y80VDD_X90Y80VSS X90Y80VDDDM X90Y80VSS 0
I_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VDDDM 0.8 AC=1
V_X90Y90VDD_X90Y90VSS X90Y90VDDDM X90Y90VSS 0
I_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VDDDM 0.8 AC=1
V_X90Y100VDD_X90Y100VSS X90Y100VDDDM X90Y100VSS 0
I_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VDDDM 0.8 AC=1
V_X90Y110VDD_X90Y110VSS X90Y110VDDDM X90Y110VSS 0
I_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VDDDM 0.8 AC=1
V_X100Y120VDD_X100Y120VSS X100Y120VDDDM X100Y120VSS 0
I_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VDDDM 0.8 AC=1
V_X100Y10VDD_X100Y10VSS X100Y10VDDDM X100Y10VSS 0
I_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VDDDM 0.8 AC=1
V_X100Y20VDD_X100Y20VSS X100Y20VDDDM X100Y20VSS 0
I_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VDDDM 0.8 AC=1
V_X100Y30VDD_X100Y30VSS X100Y30VDDDM X100Y30VSS 0
I_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VDDDM 0.8 AC=1
V_X100Y40VDD_X100Y40VSS X100Y40VDDDM X100Y40VSS 0
I_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VDDDM 0.8 AC=1
V_X100Y50VDD_X100Y50VSS X100Y50VDDDM X100Y50VSS 0
I_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VDDDM 0.8 AC=1
V_X100Y60VDD_X100Y60VSS X100Y60VDDDM X100Y60VSS 0
I_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VDDDM 0.8 AC=1
V_X100Y70VDD_X100Y70VSS X100Y70VDDDM X100Y70VSS 0
I_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VDDDM 0.8 AC=1
V_X100Y80VDD_X100Y80VSS X100Y80VDDDM X100Y80VSS 0
I_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VDDDM 0.8 AC=1
V_X100Y90VDD_X100Y90VSS X100Y90VDDDM X100Y90VSS 0
I_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VDDDM 0.8 AC=1
V_X100Y100VDD_X100Y100VSS X100Y100VDDDM X100Y100VSS 0
I_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VDDDM 0.8 AC=1
V_X100Y110VDD_X100Y110VSS X100Y110VDDDM X100Y110VSS 0
I_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VDDDM 0.8 AC=1
V_X110Y120VDD_X110Y120VSS X110Y120VDDDM X110Y120VSS 0
I_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VDDDM 0.8 AC=1
V_X110Y10VDD_X110Y10VSS X110Y10VDDDM X110Y10VSS 0
I_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VDDDM 0.8 AC=1
V_X110Y20VDD_X110Y20VSS X110Y20VDDDM X110Y20VSS 0
I_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VDDDM 0.8 AC=1
V_X110Y30VDD_X110Y30VSS X110Y30VDDDM X110Y30VSS 0
I_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VDDDM 0.8 AC=1
V_X110Y40VDD_X110Y40VSS X110Y40VDDDM X110Y40VSS 0
I_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VDDDM 0.8 AC=1
V_X110Y50VDD_X110Y50VSS X110Y50VDDDM X110Y50VSS 0
I_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VDDDM 0.8 AC=1
V_X110Y60VDD_X110Y60VSS X110Y60VDDDM X110Y60VSS 0
I_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VDDDM 0.8 AC=1
V_X110Y70VDD_X110Y70VSS X110Y70VDDDM X110Y70VSS 0
I_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VDDDM 0.8 AC=1
V_X110Y80VDD_X110Y80VSS X110Y80VDDDM X110Y80VSS 0
I_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VDDDM 0.8 AC=1
V_X110Y90VDD_X110Y90VSS X110Y90VDDDM X110Y90VSS 0
I_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VDDDM 0.8 AC=1
V_X110Y100VDD_X110Y100VSS X110Y100VDDDM X110Y100VSS 0
I_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VDDDM 0.8 AC=1
V_X110Y110VDD_X110Y110VSS X110Y110VDDDM X110Y110VSS 0
Rs1_1 VDD 11_1 0.027Ohm
Cp1_1 11_1 VSS 131.33333333333331nF
Rs2_1 11_1 12_1 0.027Ohm
Cp2_1 12_1 VSS 213.33333333333331nF
Fs_1 12_1 VSS V_X60Y60VDD_X60Y60VSS 3.0
Rg_1 VSS X60Y60VSS 0.025Ohm
Bs_1 13_1 X60Y60VSS v=(((0.3333333333333333+((v(Vref_1)-v(X60Y60VDD,X60Y60VSS))*3.0))<1?((0.3333333333333333+((v(Vref_1)-v(X60Y60VDD,X60Y60VSS))*3.0))>0?(0.3333333333333333+((v(Vref_1)-v(X60Y60VDD,X60Y60VSS))*3.0)):0):1)*v(VDD,VSS))
Rs3_1 13_1 14_1 0.009Ohm
Cp3_1 14_1 X60Y60VSS 394nF
Rs4_1 14_1 X60Y60VDD 0.009Ohm
Cp4_1 X60Y60VDD X60Y60VSS 640nF
Vref_1 Vref_1 0 1.1
.ends dut
XRegulator0 VDD0 VSS0 Regulator
Rgnd VSS0 0 0
XPcbModelLumped0 VDD0 VSS0 VDD1 VSS1 PcbModelLumped
XChipPackage1 VDD1 VSS1 VDD2 VSS2 ChipPackage
XChipBump2 VDD2 VSS2 VDD3 VSS3 ChipBump
Xdut3 VDD3 VSS3 dut


# distributed feedback
.title 20200622-105452
.option rshunt = 1.0e12
.subckt PcbBuckConverter VDD VSS
C1 VDD 12 2340uF
R1 12 13 0Ohm
L1 13 VSS 0nH
C2 VDD 22 0uF
R2 22 23 1000000000000.0Ohm
L2 23 VSS 0nH
Ls VDD 31 0.33uH
Rs 31 32 20mOhm
Vs 32 VSS 1.1
.ends PcbBuckConverter

.subckt PcbModelLumped VDD1 VSS1 VDD2 VSS2
Rs1 VDD1 11 1000mOhm
Ls1 11 VDD2 0nH
Rs2 VSS1 21 1000mOhm
Ls2 21 VSS2 0nH
Rp VDD2 VDD2M 0mOhm
Cp VDD2M VSS2 0uF
.ends PcbModelLumped

.subckt dut VDD VSS
R_X10Y10VDD_X20Y10VDD X10Y10VDD X15Y10VDD 25mOhm
L_X10Y10VDD_X20Y10VDD X15Y10VDD X20Y10VDD 2.91e-06nH
R_X10Y10VSS_X20Y10VSS X10Y10VSS X15Y10VSS 25mOhm
L_X10Y10VSS_X20Y10VSS X15Y10VSS X20Y10VSS 2.91e-06nH
R_X20Y10VDD_X30Y10VDD X20Y10VDD X25Y10VDD 25mOhm
L_X20Y10VDD_X30Y10VDD X25Y10VDD X30Y10VDD 2.91e-06nH
R_X20Y10VSS_X30Y10VSS X20Y10VSS X25Y10VSS 25mOhm
L_X20Y10VSS_X30Y10VSS X25Y10VSS X30Y10VSS 2.91e-06nH
R_X30Y10VDD_X40Y10VDD X30Y10VDD X35Y10VDD 25mOhm
L_X30Y10VDD_X40Y10VDD X35Y10VDD X40Y10VDD 2.91e-06nH
R_X30Y10VSS_X40Y10VSS X30Y10VSS X35Y10VSS 25mOhm
L_X30Y10VSS_X40Y10VSS X35Y10VSS X40Y10VSS 2.91e-06nH
R_X40Y10VDD_X50Y10VDD X40Y10VDD X45Y10VDD 25mOhm
L_X40Y10VDD_X50Y10VDD X45Y10VDD X50Y10VDD 2.91e-06nH
R_X40Y10VSS_X50Y10VSS X40Y10VSS X45Y10VSS 25mOhm
L_X40Y10VSS_X50Y10VSS X45Y10VSS X50Y10VSS 2.91e-06nH
R_X50Y10VDD_X60Y10VDD X50Y10VDD X55Y10VDD 25mOhm
L_X50Y10VDD_X60Y10VDD X55Y10VDD X60Y10VDD 2.91e-06nH
R_X50Y10VSS_X60Y10VSS X50Y10VSS X55Y10VSS 25mOhm
L_X50Y10VSS_X60Y10VSS X55Y10VSS X60Y10VSS 2.91e-06nH
R_X60Y10VDD_X70Y10VDD X60Y10VDD X65Y10VDD 25mOhm
L_X60Y10VDD_X70Y10VDD X65Y10VDD X70Y10VDD 2.91e-06nH
R_X60Y10VSS_X70Y10VSS X60Y10VSS X65Y10VSS 25mOhm
L_X60Y10VSS_X70Y10VSS X65Y10VSS X70Y10VSS 2.91e-06nH
R_X70Y10VDD_X80Y10VDD X70Y10VDD X75Y10VDD 25mOhm
L_X70Y10VDD_X80Y10VDD X75Y10VDD X80Y10VDD 2.91e-06nH
R_X70Y10VSS_X80Y10VSS X70Y10VSS X75Y10VSS 25mOhm
L_X70Y10VSS_X80Y10VSS X75Y10VSS X80Y10VSS 2.91e-06nH
R_X80Y10VDD_X90Y10VDD X80Y10VDD X85Y10VDD 25mOhm
L_X80Y10VDD_X90Y10VDD X85Y10VDD X90Y10VDD 2.91e-06nH
R_X80Y10VSS_X90Y10VSS X80Y10VSS X85Y10VSS 25mOhm
L_X80Y10VSS_X90Y10VSS X85Y10VSS X90Y10VSS 2.91e-06nH
R_X90Y10VDD_X100Y10VDD X90Y10VDD X95Y10VDD 25mOhm
L_X90Y10VDD_X100Y10VDD X95Y10VDD X100Y10VDD 2.91e-06nH
R_X90Y10VSS_X100Y10VSS X90Y10VSS X95Y10VSS 25mOhm
L_X90Y10VSS_X100Y10VSS X95Y10VSS X100Y10VSS 2.91e-06nH
R_X100Y10VDD_X110Y10VDD X100Y10VDD X105Y10VDD 25mOhm
L_X100Y10VDD_X110Y10VDD X105Y10VDD X110Y10VDD 2.91e-06nH
R_X100Y10VSS_X110Y10VSS X100Y10VSS X105Y10VSS 25mOhm
L_X100Y10VSS_X110Y10VSS X105Y10VSS X110Y10VSS 2.91e-06nH
R_X110Y10VDD_X120Y10VDD X110Y10VDD X115Y10VDD 25mOhm
L_X110Y10VDD_X120Y10VDD X115Y10VDD X120Y10VDD 2.91e-06nH
R_X110Y10VSS_X120Y10VSS X110Y10VSS X115Y10VSS 25mOhm
L_X110Y10VSS_X120Y10VSS X115Y10VSS X120Y10VSS 2.91e-06nH
R_X10Y20VDD_X20Y20VDD X10Y20VDD X15Y20VDD 25mOhm
L_X10Y20VDD_X20Y20VDD X15Y20VDD X20Y20VDD 2.91e-06nH
R_X10Y20VSS_X20Y20VSS X10Y20VSS X15Y20VSS 25mOhm
L_X10Y20VSS_X20Y20VSS X15Y20VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X30Y20VDD X20Y20VDD X25Y20VDD 25mOhm
L_X20Y20VDD_X30Y20VDD X25Y20VDD X30Y20VDD 2.91e-06nH
R_X20Y20VSS_X30Y20VSS X20Y20VSS X25Y20VSS 25mOhm
L_X20Y20VSS_X30Y20VSS X25Y20VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X40Y20VDD X30Y20VDD X35Y20VDD 25mOhm
L_X30Y20VDD_X40Y20VDD X35Y20VDD X40Y20VDD 2.91e-06nH
R_X30Y20VSS_X40Y20VSS X30Y20VSS X35Y20VSS 25mOhm
L_X30Y20VSS_X40Y20VSS X35Y20VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X50Y20VDD X40Y20VDD X45Y20VDD 25mOhm
L_X40Y20VDD_X50Y20VDD X45Y20VDD X50Y20VDD 2.91e-06nH
R_X40Y20VSS_X50Y20VSS X40Y20VSS X45Y20VSS 25mOhm
L_X40Y20VSS_X50Y20VSS X45Y20VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X60Y20VDD X50Y20VDD X55Y20VDD 25mOhm
L_X50Y20VDD_X60Y20VDD X55Y20VDD X60Y20VDD 2.91e-06nH
R_X50Y20VSS_X60Y20VSS X50Y20VSS X55Y20VSS 25mOhm
L_X50Y20VSS_X60Y20VSS X55Y20VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X70Y20VDD X60Y20VDD X65Y20VDD 25mOhm
L_X60Y20VDD_X70Y20VDD X65Y20VDD X70Y20VDD 2.91e-06nH
R_X60Y20VSS_X70Y20VSS X60Y20VSS X65Y20VSS 25mOhm
L_X60Y20VSS_X70Y20VSS X65Y20VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X80Y20VDD X70Y20VDD X75Y20VDD 25mOhm
L_X70Y20VDD_X80Y20VDD X75Y20VDD X80Y20VDD 2.91e-06nH
R_X70Y20VSS_X80Y20VSS X70Y20VSS X75Y20VSS 25mOhm
L_X70Y20VSS_X80Y20VSS X75Y20VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X90Y20VDD X80Y20VDD X85Y20VDD 25mOhm
L_X80Y20VDD_X90Y20VDD X85Y20VDD X90Y20VDD 2.91e-06nH
R_X80Y20VSS_X90Y20VSS X80Y20VSS X85Y20VSS 25mOhm
L_X80Y20VSS_X90Y20VSS X85Y20VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X100Y20VDD X90Y20VDD X95Y20VDD 25mOhm
L_X90Y20VDD_X100Y20VDD X95Y20VDD X100Y20VDD 2.91e-06nH
R_X90Y20VSS_X100Y20VSS X90Y20VSS X95Y20VSS 25mOhm
L_X90Y20VSS_X100Y20VSS X95Y20VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X110Y20VDD X100Y20VDD X105Y20VDD 25mOhm
L_X100Y20VDD_X110Y20VDD X105Y20VDD X110Y20VDD 2.91e-06nH
R_X100Y20VSS_X110Y20VSS X100Y20VSS X105Y20VSS 25mOhm
L_X100Y20VSS_X110Y20VSS X105Y20VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X120Y20VDD X110Y20VDD X115Y20VDD 25mOhm
L_X110Y20VDD_X120Y20VDD X115Y20VDD X120Y20VDD 2.91e-06nH
R_X110Y20VSS_X120Y20VSS X110Y20VSS X115Y20VSS 25mOhm
L_X110Y20VSS_X120Y20VSS X115Y20VSS X120Y20VSS 2.91e-06nH
R_X10Y30VDD_X20Y30VDD X10Y30VDD X15Y30VDD 25mOhm
L_X10Y30VDD_X20Y30VDD X15Y30VDD X20Y30VDD 2.91e-06nH
R_X10Y30VSS_X20Y30VSS X10Y30VSS X15Y30VSS 25mOhm
L_X10Y30VSS_X20Y30VSS X15Y30VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X30Y30VDD X20Y30VDD X25Y30VDD 25mOhm
L_X20Y30VDD_X30Y30VDD X25Y30VDD X30Y30VDD 2.91e-06nH
R_X20Y30VSS_X30Y30VSS X20Y30VSS X25Y30VSS 25mOhm
L_X20Y30VSS_X30Y30VSS X25Y30VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X40Y30VDD X30Y30VDD X35Y30VDD 25mOhm
L_X30Y30VDD_X40Y30VDD X35Y30VDD X40Y30VDD 2.91e-06nH
R_X30Y30VSS_X40Y30VSS X30Y30VSS X35Y30VSS 25mOhm
L_X30Y30VSS_X40Y30VSS X35Y30VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X50Y30VDD X40Y30VDD X45Y30VDD 25mOhm
L_X40Y30VDD_X50Y30VDD X45Y30VDD X50Y30VDD 2.91e-06nH
R_X40Y30VSS_X50Y30VSS X40Y30VSS X45Y30VSS 25mOhm
L_X40Y30VSS_X50Y30VSS X45Y30VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X60Y30VDD X50Y30VDD X55Y30VDD 25mOhm
L_X50Y30VDD_X60Y30VDD X55Y30VDD X60Y30VDD 2.91e-06nH
R_X50Y30VSS_X60Y30VSS X50Y30VSS X55Y30VSS 25mOhm
L_X50Y30VSS_X60Y30VSS X55Y30VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X70Y30VDD X60Y30VDD X65Y30VDD 25mOhm
L_X60Y30VDD_X70Y30VDD X65Y30VDD X70Y30VDD 2.91e-06nH
R_X60Y30VSS_X70Y30VSS X60Y30VSS X65Y30VSS 25mOhm
L_X60Y30VSS_X70Y30VSS X65Y30VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X80Y30VDD X70Y30VDD X75Y30VDD 25mOhm
L_X70Y30VDD_X80Y30VDD X75Y30VDD X80Y30VDD 2.91e-06nH
R_X70Y30VSS_X80Y30VSS X70Y30VSS X75Y30VSS 25mOhm
L_X70Y30VSS_X80Y30VSS X75Y30VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X90Y30VDD X80Y30VDD X85Y30VDD 25mOhm
L_X80Y30VDD_X90Y30VDD X85Y30VDD X90Y30VDD 2.91e-06nH
R_X80Y30VSS_X90Y30VSS X80Y30VSS X85Y30VSS 25mOhm
L_X80Y30VSS_X90Y30VSS X85Y30VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X100Y30VDD X90Y30VDD X95Y30VDD 25mOhm
L_X90Y30VDD_X100Y30VDD X95Y30VDD X100Y30VDD 2.91e-06nH
R_X90Y30VSS_X100Y30VSS X90Y30VSS X95Y30VSS 25mOhm
L_X90Y30VSS_X100Y30VSS X95Y30VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X110Y30VDD X100Y30VDD X105Y30VDD 25mOhm
L_X100Y30VDD_X110Y30VDD X105Y30VDD X110Y30VDD 2.91e-06nH
R_X100Y30VSS_X110Y30VSS X100Y30VSS X105Y30VSS 25mOhm
L_X100Y30VSS_X110Y30VSS X105Y30VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X120Y30VDD X110Y30VDD X115Y30VDD 25mOhm
L_X110Y30VDD_X120Y30VDD X115Y30VDD X120Y30VDD 2.91e-06nH
R_X110Y30VSS_X120Y30VSS X110Y30VSS X115Y30VSS 25mOhm
L_X110Y30VSS_X120Y30VSS X115Y30VSS X120Y30VSS 2.91e-06nH
R_X10Y40VDD_X20Y40VDD X10Y40VDD X15Y40VDD 25mOhm
L_X10Y40VDD_X20Y40VDD X15Y40VDD X20Y40VDD 2.91e-06nH
R_X10Y40VSS_X20Y40VSS X10Y40VSS X15Y40VSS 25mOhm
L_X10Y40VSS_X20Y40VSS X15Y40VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X30Y40VDD X20Y40VDD X25Y40VDD 25mOhm
L_X20Y40VDD_X30Y40VDD X25Y40VDD X30Y40VDD 2.91e-06nH
R_X20Y40VSS_X30Y40VSS X20Y40VSS X25Y40VSS 25mOhm
L_X20Y40VSS_X30Y40VSS X25Y40VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X40Y40VDD X30Y40VDD X35Y40VDD 25mOhm
L_X30Y40VDD_X40Y40VDD X35Y40VDD X40Y40VDD 2.91e-06nH
R_X30Y40VSS_X40Y40VSS X30Y40VSS X35Y40VSS 25mOhm
L_X30Y40VSS_X40Y40VSS X35Y40VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X50Y40VDD X40Y40VDD X45Y40VDD 25mOhm
L_X40Y40VDD_X50Y40VDD X45Y40VDD X50Y40VDD 2.91e-06nH
R_X40Y40VSS_X50Y40VSS X40Y40VSS X45Y40VSS 25mOhm
L_X40Y40VSS_X50Y40VSS X45Y40VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X60Y40VDD X50Y40VDD X55Y40VDD 25mOhm
L_X50Y40VDD_X60Y40VDD X55Y40VDD X60Y40VDD 2.91e-06nH
R_X50Y40VSS_X60Y40VSS X50Y40VSS X55Y40VSS 25mOhm
L_X50Y40VSS_X60Y40VSS X55Y40VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X70Y40VDD X60Y40VDD X65Y40VDD 25mOhm
L_X60Y40VDD_X70Y40VDD X65Y40VDD X70Y40VDD 2.91e-06nH
R_X60Y40VSS_X70Y40VSS X60Y40VSS X65Y40VSS 25mOhm
L_X60Y40VSS_X70Y40VSS X65Y40VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X80Y40VDD X70Y40VDD X75Y40VDD 25mOhm
L_X70Y40VDD_X80Y40VDD X75Y40VDD X80Y40VDD 2.91e-06nH
R_X70Y40VSS_X80Y40VSS X70Y40VSS X75Y40VSS 25mOhm
L_X70Y40VSS_X80Y40VSS X75Y40VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X90Y40VDD X80Y40VDD X85Y40VDD 25mOhm
L_X80Y40VDD_X90Y40VDD X85Y40VDD X90Y40VDD 2.91e-06nH
R_X80Y40VSS_X90Y40VSS X80Y40VSS X85Y40VSS 25mOhm
L_X80Y40VSS_X90Y40VSS X85Y40VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X100Y40VDD X90Y40VDD X95Y40VDD 25mOhm
L_X90Y40VDD_X100Y40VDD X95Y40VDD X100Y40VDD 2.91e-06nH
R_X90Y40VSS_X100Y40VSS X90Y40VSS X95Y40VSS 25mOhm
L_X90Y40VSS_X100Y40VSS X95Y40VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X110Y40VDD X100Y40VDD X105Y40VDD 25mOhm
L_X100Y40VDD_X110Y40VDD X105Y40VDD X110Y40VDD 2.91e-06nH
R_X100Y40VSS_X110Y40VSS X100Y40VSS X105Y40VSS 25mOhm
L_X100Y40VSS_X110Y40VSS X105Y40VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X120Y40VDD X110Y40VDD X115Y40VDD 25mOhm
L_X110Y40VDD_X120Y40VDD X115Y40VDD X120Y40VDD 2.91e-06nH
R_X110Y40VSS_X120Y40VSS X110Y40VSS X115Y40VSS 25mOhm
L_X110Y40VSS_X120Y40VSS X115Y40VSS X120Y40VSS 2.91e-06nH
R_X10Y50VDD_X20Y50VDD X10Y50VDD X15Y50VDD 25mOhm
L_X10Y50VDD_X20Y50VDD X15Y50VDD X20Y50VDD 2.91e-06nH
R_X10Y50VSS_X20Y50VSS X10Y50VSS X15Y50VSS 25mOhm
L_X10Y50VSS_X20Y50VSS X15Y50VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X30Y50VDD X20Y50VDD X25Y50VDD 25mOhm
L_X20Y50VDD_X30Y50VDD X25Y50VDD X30Y50VDD 2.91e-06nH
R_X20Y50VSS_X30Y50VSS X20Y50VSS X25Y50VSS 25mOhm
L_X20Y50VSS_X30Y50VSS X25Y50VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X40Y50VDD X30Y50VDD X35Y50VDD 25mOhm
L_X30Y50VDD_X40Y50VDD X35Y50VDD X40Y50VDD 2.91e-06nH
R_X30Y50VSS_X40Y50VSS X30Y50VSS X35Y50VSS 25mOhm
L_X30Y50VSS_X40Y50VSS X35Y50VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X50Y50VDD X40Y50VDD X45Y50VDD 25mOhm
L_X40Y50VDD_X50Y50VDD X45Y50VDD X50Y50VDD 2.91e-06nH
R_X40Y50VSS_X50Y50VSS X40Y50VSS X45Y50VSS 25mOhm
L_X40Y50VSS_X50Y50VSS X45Y50VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X60Y50VDD X50Y50VDD X55Y50VDD 25mOhm
L_X50Y50VDD_X60Y50VDD X55Y50VDD X60Y50VDD 2.91e-06nH
R_X50Y50VSS_X60Y50VSS X50Y50VSS X55Y50VSS 25mOhm
L_X50Y50VSS_X60Y50VSS X55Y50VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X70Y50VDD X60Y50VDD X65Y50VDD 25mOhm
L_X60Y50VDD_X70Y50VDD X65Y50VDD X70Y50VDD 2.91e-06nH
R_X60Y50VSS_X70Y50VSS X60Y50VSS X65Y50VSS 25mOhm
L_X60Y50VSS_X70Y50VSS X65Y50VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X80Y50VDD X70Y50VDD X75Y50VDD 25mOhm
L_X70Y50VDD_X80Y50VDD X75Y50VDD X80Y50VDD 2.91e-06nH
R_X70Y50VSS_X80Y50VSS X70Y50VSS X75Y50VSS 25mOhm
L_X70Y50VSS_X80Y50VSS X75Y50VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X90Y50VDD X80Y50VDD X85Y50VDD 25mOhm
L_X80Y50VDD_X90Y50VDD X85Y50VDD X90Y50VDD 2.91e-06nH
R_X80Y50VSS_X90Y50VSS X80Y50VSS X85Y50VSS 25mOhm
L_X80Y50VSS_X90Y50VSS X85Y50VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X100Y50VDD X90Y50VDD X95Y50VDD 25mOhm
L_X90Y50VDD_X100Y50VDD X95Y50VDD X100Y50VDD 2.91e-06nH
R_X90Y50VSS_X100Y50VSS X90Y50VSS X95Y50VSS 25mOhm
L_X90Y50VSS_X100Y50VSS X95Y50VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X110Y50VDD X100Y50VDD X105Y50VDD 25mOhm
L_X100Y50VDD_X110Y50VDD X105Y50VDD X110Y50VDD 2.91e-06nH
R_X100Y50VSS_X110Y50VSS X100Y50VSS X105Y50VSS 25mOhm
L_X100Y50VSS_X110Y50VSS X105Y50VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X120Y50VDD X110Y50VDD X115Y50VDD 25mOhm
L_X110Y50VDD_X120Y50VDD X115Y50VDD X120Y50VDD 2.91e-06nH
R_X110Y50VSS_X120Y50VSS X110Y50VSS X115Y50VSS 25mOhm
L_X110Y50VSS_X120Y50VSS X115Y50VSS X120Y50VSS 2.91e-06nH
R_X10Y60VDD_X20Y60VDD X10Y60VDD X15Y60VDD 25mOhm
L_X10Y60VDD_X20Y60VDD X15Y60VDD X20Y60VDD 2.91e-06nH
R_X10Y60VSS_X20Y60VSS X10Y60VSS X15Y60VSS 25mOhm
L_X10Y60VSS_X20Y60VSS X15Y60VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X30Y60VDD X20Y60VDD X25Y60VDD 25mOhm
L_X20Y60VDD_X30Y60VDD X25Y60VDD X30Y60VDD 2.91e-06nH
R_X20Y60VSS_X30Y60VSS X20Y60VSS X25Y60VSS 25mOhm
L_X20Y60VSS_X30Y60VSS X25Y60VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X40Y60VDD X30Y60VDD X35Y60VDD 25mOhm
L_X30Y60VDD_X40Y60VDD X35Y60VDD X40Y60VDD 2.91e-06nH
R_X30Y60VSS_X40Y60VSS X30Y60VSS X35Y60VSS 25mOhm
L_X30Y60VSS_X40Y60VSS X35Y60VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X50Y60VDD X40Y60VDD X45Y60VDD 25mOhm
L_X40Y60VDD_X50Y60VDD X45Y60VDD X50Y60VDD 2.91e-06nH
R_X40Y60VSS_X50Y60VSS X40Y60VSS X45Y60VSS 25mOhm
L_X40Y60VSS_X50Y60VSS X45Y60VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X60Y60VDD X50Y60VDD X55Y60VDD 25mOhm
L_X50Y60VDD_X60Y60VDD X55Y60VDD X60Y60VDD 2.91e-06nH
R_X50Y60VSS_X60Y60VSS X50Y60VSS X55Y60VSS 25mOhm
L_X50Y60VSS_X60Y60VSS X55Y60VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X70Y60VDD X60Y60VDD X65Y60VDD 25mOhm
L_X60Y60VDD_X70Y60VDD X65Y60VDD X70Y60VDD 2.91e-06nH
R_X60Y60VSS_X70Y60VSS X60Y60VSS X65Y60VSS 25mOhm
L_X60Y60VSS_X70Y60VSS X65Y60VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X80Y60VDD X70Y60VDD X75Y60VDD 25mOhm
L_X70Y60VDD_X80Y60VDD X75Y60VDD X80Y60VDD 2.91e-06nH
R_X70Y60VSS_X80Y60VSS X70Y60VSS X75Y60VSS 25mOhm
L_X70Y60VSS_X80Y60VSS X75Y60VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X90Y60VDD X80Y60VDD X85Y60VDD 25mOhm
L_X80Y60VDD_X90Y60VDD X85Y60VDD X90Y60VDD 2.91e-06nH
R_X80Y60VSS_X90Y60VSS X80Y60VSS X85Y60VSS 25mOhm
L_X80Y60VSS_X90Y60VSS X85Y60VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X100Y60VDD X90Y60VDD X95Y60VDD 25mOhm
L_X90Y60VDD_X100Y60VDD X95Y60VDD X100Y60VDD 2.91e-06nH
R_X90Y60VSS_X100Y60VSS X90Y60VSS X95Y60VSS 25mOhm
L_X90Y60VSS_X100Y60VSS X95Y60VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X110Y60VDD X100Y60VDD X105Y60VDD 25mOhm
L_X100Y60VDD_X110Y60VDD X105Y60VDD X110Y60VDD 2.91e-06nH
R_X100Y60VSS_X110Y60VSS X100Y60VSS X105Y60VSS 25mOhm
L_X100Y60VSS_X110Y60VSS X105Y60VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X120Y60VDD X110Y60VDD X115Y60VDD 25mOhm
L_X110Y60VDD_X120Y60VDD X115Y60VDD X120Y60VDD 2.91e-06nH
R_X110Y60VSS_X120Y60VSS X110Y60VSS X115Y60VSS 25mOhm
L_X110Y60VSS_X120Y60VSS X115Y60VSS X120Y60VSS 2.91e-06nH
R_X10Y70VDD_X20Y70VDD X10Y70VDD X15Y70VDD 25mOhm
L_X10Y70VDD_X20Y70VDD X15Y70VDD X20Y70VDD 2.91e-06nH
R_X10Y70VSS_X20Y70VSS X10Y70VSS X15Y70VSS 25mOhm
L_X10Y70VSS_X20Y70VSS X15Y70VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X30Y70VDD X20Y70VDD X25Y70VDD 25mOhm
L_X20Y70VDD_X30Y70VDD X25Y70VDD X30Y70VDD 2.91e-06nH
R_X20Y70VSS_X30Y70VSS X20Y70VSS X25Y70VSS 25mOhm
L_X20Y70VSS_X30Y70VSS X25Y70VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X40Y70VDD X30Y70VDD X35Y70VDD 25mOhm
L_X30Y70VDD_X40Y70VDD X35Y70VDD X40Y70VDD 2.91e-06nH
R_X30Y70VSS_X40Y70VSS X30Y70VSS X35Y70VSS 25mOhm
L_X30Y70VSS_X40Y70VSS X35Y70VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X50Y70VDD X40Y70VDD X45Y70VDD 25mOhm
L_X40Y70VDD_X50Y70VDD X45Y70VDD X50Y70VDD 2.91e-06nH
R_X40Y70VSS_X50Y70VSS X40Y70VSS X45Y70VSS 25mOhm
L_X40Y70VSS_X50Y70VSS X45Y70VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X60Y70VDD X50Y70VDD X55Y70VDD 25mOhm
L_X50Y70VDD_X60Y70VDD X55Y70VDD X60Y70VDD 2.91e-06nH
R_X50Y70VSS_X60Y70VSS X50Y70VSS X55Y70VSS 25mOhm
L_X50Y70VSS_X60Y70VSS X55Y70VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X70Y70VDD X60Y70VDD X65Y70VDD 25mOhm
L_X60Y70VDD_X70Y70VDD X65Y70VDD X70Y70VDD 2.91e-06nH
R_X60Y70VSS_X70Y70VSS X60Y70VSS X65Y70VSS 25mOhm
L_X60Y70VSS_X70Y70VSS X65Y70VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X80Y70VDD X70Y70VDD X75Y70VDD 25mOhm
L_X70Y70VDD_X80Y70VDD X75Y70VDD X80Y70VDD 2.91e-06nH
R_X70Y70VSS_X80Y70VSS X70Y70VSS X75Y70VSS 25mOhm
L_X70Y70VSS_X80Y70VSS X75Y70VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X90Y70VDD X80Y70VDD X85Y70VDD 25mOhm
L_X80Y70VDD_X90Y70VDD X85Y70VDD X90Y70VDD 2.91e-06nH
R_X80Y70VSS_X90Y70VSS X80Y70VSS X85Y70VSS 25mOhm
L_X80Y70VSS_X90Y70VSS X85Y70VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X100Y70VDD X90Y70VDD X95Y70VDD 25mOhm
L_X90Y70VDD_X100Y70VDD X95Y70VDD X100Y70VDD 2.91e-06nH
R_X90Y70VSS_X100Y70VSS X90Y70VSS X95Y70VSS 25mOhm
L_X90Y70VSS_X100Y70VSS X95Y70VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X110Y70VDD X100Y70VDD X105Y70VDD 25mOhm
L_X100Y70VDD_X110Y70VDD X105Y70VDD X110Y70VDD 2.91e-06nH
R_X100Y70VSS_X110Y70VSS X100Y70VSS X105Y70VSS 25mOhm
L_X100Y70VSS_X110Y70VSS X105Y70VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X120Y70VDD X110Y70VDD X115Y70VDD 25mOhm
L_X110Y70VDD_X120Y70VDD X115Y70VDD X120Y70VDD 2.91e-06nH
R_X110Y70VSS_X120Y70VSS X110Y70VSS X115Y70VSS 25mOhm
L_X110Y70VSS_X120Y70VSS X115Y70VSS X120Y70VSS 2.91e-06nH
R_X10Y80VDD_X20Y80VDD X10Y80VDD X15Y80VDD 25mOhm
L_X10Y80VDD_X20Y80VDD X15Y80VDD X20Y80VDD 2.91e-06nH
R_X10Y80VSS_X20Y80VSS X10Y80VSS X15Y80VSS 25mOhm
L_X10Y80VSS_X20Y80VSS X15Y80VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X30Y80VDD X20Y80VDD X25Y80VDD 25mOhm
L_X20Y80VDD_X30Y80VDD X25Y80VDD X30Y80VDD 2.91e-06nH
R_X20Y80VSS_X30Y80VSS X20Y80VSS X25Y80VSS 25mOhm
L_X20Y80VSS_X30Y80VSS X25Y80VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X40Y80VDD X30Y80VDD X35Y80VDD 25mOhm
L_X30Y80VDD_X40Y80VDD X35Y80VDD X40Y80VDD 2.91e-06nH
R_X30Y80VSS_X40Y80VSS X30Y80VSS X35Y80VSS 25mOhm
L_X30Y80VSS_X40Y80VSS X35Y80VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X50Y80VDD X40Y80VDD X45Y80VDD 25mOhm
L_X40Y80VDD_X50Y80VDD X45Y80VDD X50Y80VDD 2.91e-06nH
R_X40Y80VSS_X50Y80VSS X40Y80VSS X45Y80VSS 25mOhm
L_X40Y80VSS_X50Y80VSS X45Y80VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X60Y80VDD X50Y80VDD X55Y80VDD 25mOhm
L_X50Y80VDD_X60Y80VDD X55Y80VDD X60Y80VDD 2.91e-06nH
R_X50Y80VSS_X60Y80VSS X50Y80VSS X55Y80VSS 25mOhm
L_X50Y80VSS_X60Y80VSS X55Y80VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X70Y80VDD X60Y80VDD X65Y80VDD 25mOhm
L_X60Y80VDD_X70Y80VDD X65Y80VDD X70Y80VDD 2.91e-06nH
R_X60Y80VSS_X70Y80VSS X60Y80VSS X65Y80VSS 25mOhm
L_X60Y80VSS_X70Y80VSS X65Y80VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X80Y80VDD X70Y80VDD X75Y80VDD 25mOhm
L_X70Y80VDD_X80Y80VDD X75Y80VDD X80Y80VDD 2.91e-06nH
R_X70Y80VSS_X80Y80VSS X70Y80VSS X75Y80VSS 25mOhm
L_X70Y80VSS_X80Y80VSS X75Y80VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X90Y80VDD X80Y80VDD X85Y80VDD 25mOhm
L_X80Y80VDD_X90Y80VDD X85Y80VDD X90Y80VDD 2.91e-06nH
R_X80Y80VSS_X90Y80VSS X80Y80VSS X85Y80VSS 25mOhm
L_X80Y80VSS_X90Y80VSS X85Y80VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X100Y80VDD X90Y80VDD X95Y80VDD 25mOhm
L_X90Y80VDD_X100Y80VDD X95Y80VDD X100Y80VDD 2.91e-06nH
R_X90Y80VSS_X100Y80VSS X90Y80VSS X95Y80VSS 25mOhm
L_X90Y80VSS_X100Y80VSS X95Y80VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X110Y80VDD X100Y80VDD X105Y80VDD 25mOhm
L_X100Y80VDD_X110Y80VDD X105Y80VDD X110Y80VDD 2.91e-06nH
R_X100Y80VSS_X110Y80VSS X100Y80VSS X105Y80VSS 25mOhm
L_X100Y80VSS_X110Y80VSS X105Y80VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X120Y80VDD X110Y80VDD X115Y80VDD 25mOhm
L_X110Y80VDD_X120Y80VDD X115Y80VDD X120Y80VDD 2.91e-06nH
R_X110Y80VSS_X120Y80VSS X110Y80VSS X115Y80VSS 25mOhm
L_X110Y80VSS_X120Y80VSS X115Y80VSS X120Y80VSS 2.91e-06nH
R_X10Y90VDD_X20Y90VDD X10Y90VDD X15Y90VDD 25mOhm
L_X10Y90VDD_X20Y90VDD X15Y90VDD X20Y90VDD 2.91e-06nH
R_X10Y90VSS_X20Y90VSS X10Y90VSS X15Y90VSS 25mOhm
L_X10Y90VSS_X20Y90VSS X15Y90VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X30Y90VDD X20Y90VDD X25Y90VDD 25mOhm
L_X20Y90VDD_X30Y90VDD X25Y90VDD X30Y90VDD 2.91e-06nH
R_X20Y90VSS_X30Y90VSS X20Y90VSS X25Y90VSS 25mOhm
L_X20Y90VSS_X30Y90VSS X25Y90VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X40Y90VDD X30Y90VDD X35Y90VDD 25mOhm
L_X30Y90VDD_X40Y90VDD X35Y90VDD X40Y90VDD 2.91e-06nH
R_X30Y90VSS_X40Y90VSS X30Y90VSS X35Y90VSS 25mOhm
L_X30Y90VSS_X40Y90VSS X35Y90VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X50Y90VDD X40Y90VDD X45Y90VDD 25mOhm
L_X40Y90VDD_X50Y90VDD X45Y90VDD X50Y90VDD 2.91e-06nH
R_X40Y90VSS_X50Y90VSS X40Y90VSS X45Y90VSS 25mOhm
L_X40Y90VSS_X50Y90VSS X45Y90VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X60Y90VDD X50Y90VDD X55Y90VDD 25mOhm
L_X50Y90VDD_X60Y90VDD X55Y90VDD X60Y90VDD 2.91e-06nH
R_X50Y90VSS_X60Y90VSS X50Y90VSS X55Y90VSS 25mOhm
L_X50Y90VSS_X60Y90VSS X55Y90VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X70Y90VDD X60Y90VDD X65Y90VDD 25mOhm
L_X60Y90VDD_X70Y90VDD X65Y90VDD X70Y90VDD 2.91e-06nH
R_X60Y90VSS_X70Y90VSS X60Y90VSS X65Y90VSS 25mOhm
L_X60Y90VSS_X70Y90VSS X65Y90VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X80Y90VDD X70Y90VDD X75Y90VDD 25mOhm
L_X70Y90VDD_X80Y90VDD X75Y90VDD X80Y90VDD 2.91e-06nH
R_X70Y90VSS_X80Y90VSS X70Y90VSS X75Y90VSS 25mOhm
L_X70Y90VSS_X80Y90VSS X75Y90VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X90Y90VDD X80Y90VDD X85Y90VDD 25mOhm
L_X80Y90VDD_X90Y90VDD X85Y90VDD X90Y90VDD 2.91e-06nH
R_X80Y90VSS_X90Y90VSS X80Y90VSS X85Y90VSS 25mOhm
L_X80Y90VSS_X90Y90VSS X85Y90VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X100Y90VDD X90Y90VDD X95Y90VDD 25mOhm
L_X90Y90VDD_X100Y90VDD X95Y90VDD X100Y90VDD 2.91e-06nH
R_X90Y90VSS_X100Y90VSS X90Y90VSS X95Y90VSS 25mOhm
L_X90Y90VSS_X100Y90VSS X95Y90VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X110Y90VDD X100Y90VDD X105Y90VDD 25mOhm
L_X100Y90VDD_X110Y90VDD X105Y90VDD X110Y90VDD 2.91e-06nH
R_X100Y90VSS_X110Y90VSS X100Y90VSS X105Y90VSS 25mOhm
L_X100Y90VSS_X110Y90VSS X105Y90VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X120Y90VDD X110Y90VDD X115Y90VDD 25mOhm
L_X110Y90VDD_X120Y90VDD X115Y90VDD X120Y90VDD 2.91e-06nH
R_X110Y90VSS_X120Y90VSS X110Y90VSS X115Y90VSS 25mOhm
L_X110Y90VSS_X120Y90VSS X115Y90VSS X120Y90VSS 2.91e-06nH
R_X10Y100VDD_X20Y100VDD X10Y100VDD X15Y100VDD 25mOhm
L_X10Y100VDD_X20Y100VDD X15Y100VDD X20Y100VDD 2.91e-06nH
R_X10Y100VSS_X20Y100VSS X10Y100VSS X15Y100VSS 25mOhm
L_X10Y100VSS_X20Y100VSS X15Y100VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X30Y100VDD X20Y100VDD X25Y100VDD 25mOhm
L_X20Y100VDD_X30Y100VDD X25Y100VDD X30Y100VDD 2.91e-06nH
R_X20Y100VSS_X30Y100VSS X20Y100VSS X25Y100VSS 25mOhm
L_X20Y100VSS_X30Y100VSS X25Y100VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X40Y100VDD X30Y100VDD X35Y100VDD 25mOhm
L_X30Y100VDD_X40Y100VDD X35Y100VDD X40Y100VDD 2.91e-06nH
R_X30Y100VSS_X40Y100VSS X30Y100VSS X35Y100VSS 25mOhm
L_X30Y100VSS_X40Y100VSS X35Y100VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X50Y100VDD X40Y100VDD X45Y100VDD 25mOhm
L_X40Y100VDD_X50Y100VDD X45Y100VDD X50Y100VDD 2.91e-06nH
R_X40Y100VSS_X50Y100VSS X40Y100VSS X45Y100VSS 25mOhm
L_X40Y100VSS_X50Y100VSS X45Y100VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X60Y100VDD X50Y100VDD X55Y100VDD 25mOhm
L_X50Y100VDD_X60Y100VDD X55Y100VDD X60Y100VDD 2.91e-06nH
R_X50Y100VSS_X60Y100VSS X50Y100VSS X55Y100VSS 25mOhm
L_X50Y100VSS_X60Y100VSS X55Y100VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X70Y100VDD X60Y100VDD X65Y100VDD 25mOhm
L_X60Y100VDD_X70Y100VDD X65Y100VDD X70Y100VDD 2.91e-06nH
R_X60Y100VSS_X70Y100VSS X60Y100VSS X65Y100VSS 25mOhm
L_X60Y100VSS_X70Y100VSS X65Y100VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X80Y100VDD X70Y100VDD X75Y100VDD 25mOhm
L_X70Y100VDD_X80Y100VDD X75Y100VDD X80Y100VDD 2.91e-06nH
R_X70Y100VSS_X80Y100VSS X70Y100VSS X75Y100VSS 25mOhm
L_X70Y100VSS_X80Y100VSS X75Y100VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X90Y100VDD X80Y100VDD X85Y100VDD 25mOhm
L_X80Y100VDD_X90Y100VDD X85Y100VDD X90Y100VDD 2.91e-06nH
R_X80Y100VSS_X90Y100VSS X80Y100VSS X85Y100VSS 25mOhm
L_X80Y100VSS_X90Y100VSS X85Y100VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X100Y100VDD X90Y100VDD X95Y100VDD 25mOhm
L_X90Y100VDD_X100Y100VDD X95Y100VDD X100Y100VDD 2.91e-06nH
R_X90Y100VSS_X100Y100VSS X90Y100VSS X95Y100VSS 25mOhm
L_X90Y100VSS_X100Y100VSS X95Y100VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X110Y100VDD X100Y100VDD X105Y100VDD 25mOhm
L_X100Y100VDD_X110Y100VDD X105Y100VDD X110Y100VDD 2.91e-06nH
R_X100Y100VSS_X110Y100VSS X100Y100VSS X105Y100VSS 25mOhm
L_X100Y100VSS_X110Y100VSS X105Y100VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X120Y100VDD X110Y100VDD X115Y100VDD 25mOhm
L_X110Y100VDD_X120Y100VDD X115Y100VDD X120Y100VDD 2.91e-06nH
R_X110Y100VSS_X120Y100VSS X110Y100VSS X115Y100VSS 25mOhm
L_X110Y100VSS_X120Y100VSS X115Y100VSS X120Y100VSS 2.91e-06nH
R_X10Y110VDD_X20Y110VDD X10Y110VDD X15Y110VDD 25mOhm
L_X10Y110VDD_X20Y110VDD X15Y110VDD X20Y110VDD 2.91e-06nH
R_X10Y110VSS_X20Y110VSS X10Y110VSS X15Y110VSS 25mOhm
L_X10Y110VSS_X20Y110VSS X15Y110VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X30Y110VDD X20Y110VDD X25Y110VDD 25mOhm
L_X20Y110VDD_X30Y110VDD X25Y110VDD X30Y110VDD 2.91e-06nH
R_X20Y110VSS_X30Y110VSS X20Y110VSS X25Y110VSS 25mOhm
L_X20Y110VSS_X30Y110VSS X25Y110VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X40Y110VDD X30Y110VDD X35Y110VDD 25mOhm
L_X30Y110VDD_X40Y110VDD X35Y110VDD X40Y110VDD 2.91e-06nH
R_X30Y110VSS_X40Y110VSS X30Y110VSS X35Y110VSS 25mOhm
L_X30Y110VSS_X40Y110VSS X35Y110VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X50Y110VDD X40Y110VDD X45Y110VDD 25mOhm
L_X40Y110VDD_X50Y110VDD X45Y110VDD X50Y110VDD 2.91e-06nH
R_X40Y110VSS_X50Y110VSS X40Y110VSS X45Y110VSS 25mOhm
L_X40Y110VSS_X50Y110VSS X45Y110VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X60Y110VDD X50Y110VDD X55Y110VDD 25mOhm
L_X50Y110VDD_X60Y110VDD X55Y110VDD X60Y110VDD 2.91e-06nH
R_X50Y110VSS_X60Y110VSS X50Y110VSS X55Y110VSS 25mOhm
L_X50Y110VSS_X60Y110VSS X55Y110VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X70Y110VDD X60Y110VDD X65Y110VDD 25mOhm
L_X60Y110VDD_X70Y110VDD X65Y110VDD X70Y110VDD 2.91e-06nH
R_X60Y110VSS_X70Y110VSS X60Y110VSS X65Y110VSS 25mOhm
L_X60Y110VSS_X70Y110VSS X65Y110VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X80Y110VDD X70Y110VDD X75Y110VDD 25mOhm
L_X70Y110VDD_X80Y110VDD X75Y110VDD X80Y110VDD 2.91e-06nH
R_X70Y110VSS_X80Y110VSS X70Y110VSS X75Y110VSS 25mOhm
L_X70Y110VSS_X80Y110VSS X75Y110VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X90Y110VDD X80Y110VDD X85Y110VDD 25mOhm
L_X80Y110VDD_X90Y110VDD X85Y110VDD X90Y110VDD 2.91e-06nH
R_X80Y110VSS_X90Y110VSS X80Y110VSS X85Y110VSS 25mOhm
L_X80Y110VSS_X90Y110VSS X85Y110VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X100Y110VDD X90Y110VDD X95Y110VDD 25mOhm
L_X90Y110VDD_X100Y110VDD X95Y110VDD X100Y110VDD 2.91e-06nH
R_X90Y110VSS_X100Y110VSS X90Y110VSS X95Y110VSS 25mOhm
L_X90Y110VSS_X100Y110VSS X95Y110VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X110Y110VDD X100Y110VDD X105Y110VDD 25mOhm
L_X100Y110VDD_X110Y110VDD X105Y110VDD X110Y110VDD 2.91e-06nH
R_X100Y110VSS_X110Y110VSS X100Y110VSS X105Y110VSS 25mOhm
L_X100Y110VSS_X110Y110VSS X105Y110VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X120Y110VDD X110Y110VDD X115Y110VDD 25mOhm
L_X110Y110VDD_X120Y110VDD X115Y110VDD X120Y110VDD 2.91e-06nH
R_X110Y110VSS_X120Y110VSS X110Y110VSS X115Y110VSS 25mOhm
L_X110Y110VSS_X120Y110VSS X115Y110VSS X120Y110VSS 2.91e-06nH
R_X10Y120VDD_X20Y120VDD X10Y120VDD X15Y120VDD 25mOhm
L_X10Y120VDD_X20Y120VDD X15Y120VDD X20Y120VDD 2.91e-06nH
R_X10Y120VSS_X20Y120VSS X10Y120VSS X15Y120VSS 25mOhm
L_X10Y120VSS_X20Y120VSS X15Y120VSS X20Y120VSS 2.91e-06nH
R_X20Y120VDD_X30Y120VDD X20Y120VDD X25Y120VDD 25mOhm
L_X20Y120VDD_X30Y120VDD X25Y120VDD X30Y120VDD 2.91e-06nH
R_X20Y120VSS_X30Y120VSS X20Y120VSS X25Y120VSS 25mOhm
L_X20Y120VSS_X30Y120VSS X25Y120VSS X30Y120VSS 2.91e-06nH
R_X30Y120VDD_X40Y120VDD X30Y120VDD X35Y120VDD 25mOhm
L_X30Y120VDD_X40Y120VDD X35Y120VDD X40Y120VDD 2.91e-06nH
R_X30Y120VSS_X40Y120VSS X30Y120VSS X35Y120VSS 25mOhm
L_X30Y120VSS_X40Y120VSS X35Y120VSS X40Y120VSS 2.91e-06nH
R_X40Y120VDD_X50Y120VDD X40Y120VDD X45Y120VDD 25mOhm
L_X40Y120VDD_X50Y120VDD X45Y120VDD X50Y120VDD 2.91e-06nH
R_X40Y120VSS_X50Y120VSS X40Y120VSS X45Y120VSS 25mOhm
L_X40Y120VSS_X50Y120VSS X45Y120VSS X50Y120VSS 2.91e-06nH
R_X50Y120VDD_X60Y120VDD X50Y120VDD X55Y120VDD 25mOhm
L_X50Y120VDD_X60Y120VDD X55Y120VDD X60Y120VDD 2.91e-06nH
R_X50Y120VSS_X60Y120VSS X50Y120VSS X55Y120VSS 25mOhm
L_X50Y120VSS_X60Y120VSS X55Y120VSS X60Y120VSS 2.91e-06nH
R_X60Y120VDD_X70Y120VDD X60Y120VDD X65Y120VDD 25mOhm
L_X60Y120VDD_X70Y120VDD X65Y120VDD X70Y120VDD 2.91e-06nH
R_X60Y120VSS_X70Y120VSS X60Y120VSS X65Y120VSS 25mOhm
L_X60Y120VSS_X70Y120VSS X65Y120VSS X70Y120VSS 2.91e-06nH
R_X70Y120VDD_X80Y120VDD X70Y120VDD X75Y120VDD 25mOhm
L_X70Y120VDD_X80Y120VDD X75Y120VDD X80Y120VDD 2.91e-06nH
R_X70Y120VSS_X80Y120VSS X70Y120VSS X75Y120VSS 25mOhm
L_X70Y120VSS_X80Y120VSS X75Y120VSS X80Y120VSS 2.91e-06nH
R_X80Y120VDD_X90Y120VDD X80Y120VDD X85Y120VDD 25mOhm
L_X80Y120VDD_X90Y120VDD X85Y120VDD X90Y120VDD 2.91e-06nH
R_X80Y120VSS_X90Y120VSS X80Y120VSS X85Y120VSS 25mOhm
L_X80Y120VSS_X90Y120VSS X85Y120VSS X90Y120VSS 2.91e-06nH
R_X90Y120VDD_X100Y120VDD X90Y120VDD X95Y120VDD 25mOhm
L_X90Y120VDD_X100Y120VDD X95Y120VDD X100Y120VDD 2.91e-06nH
R_X90Y120VSS_X100Y120VSS X90Y120VSS X95Y120VSS 25mOhm
L_X90Y120VSS_X100Y120VSS X95Y120VSS X100Y120VSS 2.91e-06nH
R_X100Y120VDD_X110Y120VDD X100Y120VDD X105Y120VDD 25mOhm
L_X100Y120VDD_X110Y120VDD X105Y120VDD X110Y120VDD 2.91e-06nH
R_X100Y120VSS_X110Y120VSS X100Y120VSS X105Y120VSS 25mOhm
L_X100Y120VSS_X110Y120VSS X105Y120VSS X110Y120VSS 2.91e-06nH
R_X110Y120VDD_X120Y120VDD X110Y120VDD X115Y120VDD 25mOhm
L_X110Y120VDD_X120Y120VDD X115Y120VDD X120Y120VDD 2.91e-06nH
R_X110Y120VSS_X120Y120VSS X110Y120VSS X115Y120VSS 25mOhm
L_X110Y120VSS_X120Y120VSS X115Y120VSS X120Y120VSS 2.91e-06nH
R_X10Y10VDD_X10Y20VDD X10Y10VDD X10Y15VDD 25mOhm
L_X10Y10VDD_X10Y20VDD X10Y15VDD X10Y20VDD 2.91e-06nH
R_X10Y10VSS_X10Y20VSS X10Y10VSS X10Y15VSS 25mOhm
L_X10Y10VSS_X10Y20VSS X10Y15VSS X10Y20VSS 2.91e-06nH
R_X10Y20VDD_X10Y30VDD X10Y20VDD X10Y25VDD 25mOhm
L_X10Y20VDD_X10Y30VDD X10Y25VDD X10Y30VDD 2.91e-06nH
R_X10Y20VSS_X10Y30VSS X10Y20VSS X10Y25VSS 25mOhm
L_X10Y20VSS_X10Y30VSS X10Y25VSS X10Y30VSS 2.91e-06nH
R_X10Y30VDD_X10Y40VDD X10Y30VDD X10Y35VDD 25mOhm
L_X10Y30VDD_X10Y40VDD X10Y35VDD X10Y40VDD 2.91e-06nH
R_X10Y30VSS_X10Y40VSS X10Y30VSS X10Y35VSS 25mOhm
L_X10Y30VSS_X10Y40VSS X10Y35VSS X10Y40VSS 2.91e-06nH
R_X10Y40VDD_X10Y50VDD X10Y40VDD X10Y45VDD 25mOhm
L_X10Y40VDD_X10Y50VDD X10Y45VDD X10Y50VDD 2.91e-06nH
R_X10Y40VSS_X10Y50VSS X10Y40VSS X10Y45VSS 25mOhm
L_X10Y40VSS_X10Y50VSS X10Y45VSS X10Y50VSS 2.91e-06nH
R_X10Y50VDD_X10Y60VDD X10Y50VDD X10Y55VDD 25mOhm
L_X10Y50VDD_X10Y60VDD X10Y55VDD X10Y60VDD 2.91e-06nH
R_X10Y50VSS_X10Y60VSS X10Y50VSS X10Y55VSS 25mOhm
L_X10Y50VSS_X10Y60VSS X10Y55VSS X10Y60VSS 2.91e-06nH
R_X10Y60VDD_X10Y70VDD X10Y60VDD X10Y65VDD 25mOhm
L_X10Y60VDD_X10Y70VDD X10Y65VDD X10Y70VDD 2.91e-06nH
R_X10Y60VSS_X10Y70VSS X10Y60VSS X10Y65VSS 25mOhm
L_X10Y60VSS_X10Y70VSS X10Y65VSS X10Y70VSS 2.91e-06nH
R_X10Y70VDD_X10Y80VDD X10Y70VDD X10Y75VDD 25mOhm
L_X10Y70VDD_X10Y80VDD X10Y75VDD X10Y80VDD 2.91e-06nH
R_X10Y70VSS_X10Y80VSS X10Y70VSS X10Y75VSS 25mOhm
L_X10Y70VSS_X10Y80VSS X10Y75VSS X10Y80VSS 2.91e-06nH
R_X10Y80VDD_X10Y90VDD X10Y80VDD X10Y85VDD 25mOhm
L_X10Y80VDD_X10Y90VDD X10Y85VDD X10Y90VDD 2.91e-06nH
R_X10Y80VSS_X10Y90VSS X10Y80VSS X10Y85VSS 25mOhm
L_X10Y80VSS_X10Y90VSS X10Y85VSS X10Y90VSS 2.91e-06nH
R_X10Y90VDD_X10Y100VDD X10Y90VDD X10Y95VDD 25mOhm
L_X10Y90VDD_X10Y100VDD X10Y95VDD X10Y100VDD 2.91e-06nH
R_X10Y90VSS_X10Y100VSS X10Y90VSS X10Y95VSS 25mOhm
L_X10Y90VSS_X10Y100VSS X10Y95VSS X10Y100VSS 2.91e-06nH
R_X10Y100VDD_X10Y110VDD X10Y100VDD X10Y105VDD 25mOhm
L_X10Y100VDD_X10Y110VDD X10Y105VDD X10Y110VDD 2.91e-06nH
R_X10Y100VSS_X10Y110VSS X10Y100VSS X10Y105VSS 25mOhm
L_X10Y100VSS_X10Y110VSS X10Y105VSS X10Y110VSS 2.91e-06nH
R_X10Y110VDD_X10Y120VDD X10Y110VDD X10Y115VDD 25mOhm
L_X10Y110VDD_X10Y120VDD X10Y115VDD X10Y120VDD 2.91e-06nH
R_X10Y110VSS_X10Y120VSS X10Y110VSS X10Y115VSS 25mOhm
L_X10Y110VSS_X10Y120VSS X10Y115VSS X10Y120VSS 2.91e-06nH
R_X20Y10VDD_X20Y20VDD X20Y10VDD X20Y15VDD 25mOhm
L_X20Y10VDD_X20Y20VDD X20Y15VDD X20Y20VDD 2.91e-06nH
R_X20Y10VSS_X20Y20VSS X20Y10VSS X20Y15VSS 25mOhm
L_X20Y10VSS_X20Y20VSS X20Y15VSS X20Y20VSS 2.91e-06nH
R_X20Y20VDD_X20Y30VDD X20Y20VDD X20Y25VDD 25mOhm
L_X20Y20VDD_X20Y30VDD X20Y25VDD X20Y30VDD 2.91e-06nH
R_X20Y20VSS_X20Y30VSS X20Y20VSS X20Y25VSS 25mOhm
L_X20Y20VSS_X20Y30VSS X20Y25VSS X20Y30VSS 2.91e-06nH
R_X20Y30VDD_X20Y40VDD X20Y30VDD X20Y35VDD 25mOhm
L_X20Y30VDD_X20Y40VDD X20Y35VDD X20Y40VDD 2.91e-06nH
R_X20Y30VSS_X20Y40VSS X20Y30VSS X20Y35VSS 25mOhm
L_X20Y30VSS_X20Y40VSS X20Y35VSS X20Y40VSS 2.91e-06nH
R_X20Y40VDD_X20Y50VDD X20Y40VDD X20Y45VDD 25mOhm
L_X20Y40VDD_X20Y50VDD X20Y45VDD X20Y50VDD 2.91e-06nH
R_X20Y40VSS_X20Y50VSS X20Y40VSS X20Y45VSS 25mOhm
L_X20Y40VSS_X20Y50VSS X20Y45VSS X20Y50VSS 2.91e-06nH
R_X20Y50VDD_X20Y60VDD X20Y50VDD X20Y55VDD 25mOhm
L_X20Y50VDD_X20Y60VDD X20Y55VDD X20Y60VDD 2.91e-06nH
R_X20Y50VSS_X20Y60VSS X20Y50VSS X20Y55VSS 25mOhm
L_X20Y50VSS_X20Y60VSS X20Y55VSS X20Y60VSS 2.91e-06nH
R_X20Y60VDD_X20Y70VDD X20Y60VDD X20Y65VDD 25mOhm
L_X20Y60VDD_X20Y70VDD X20Y65VDD X20Y70VDD 2.91e-06nH
R_X20Y60VSS_X20Y70VSS X20Y60VSS X20Y65VSS 25mOhm
L_X20Y60VSS_X20Y70VSS X20Y65VSS X20Y70VSS 2.91e-06nH
R_X20Y70VDD_X20Y80VDD X20Y70VDD X20Y75VDD 25mOhm
L_X20Y70VDD_X20Y80VDD X20Y75VDD X20Y80VDD 2.91e-06nH
R_X20Y70VSS_X20Y80VSS X20Y70VSS X20Y75VSS 25mOhm
L_X20Y70VSS_X20Y80VSS X20Y75VSS X20Y80VSS 2.91e-06nH
R_X20Y80VDD_X20Y90VDD X20Y80VDD X20Y85VDD 25mOhm
L_X20Y80VDD_X20Y90VDD X20Y85VDD X20Y90VDD 2.91e-06nH
R_X20Y80VSS_X20Y90VSS X20Y80VSS X20Y85VSS 25mOhm
L_X20Y80VSS_X20Y90VSS X20Y85VSS X20Y90VSS 2.91e-06nH
R_X20Y90VDD_X20Y100VDD X20Y90VDD X20Y95VDD 25mOhm
L_X20Y90VDD_X20Y100VDD X20Y95VDD X20Y100VDD 2.91e-06nH
R_X20Y90VSS_X20Y100VSS X20Y90VSS X20Y95VSS 25mOhm
L_X20Y90VSS_X20Y100VSS X20Y95VSS X20Y100VSS 2.91e-06nH
R_X20Y100VDD_X20Y110VDD X20Y100VDD X20Y105VDD 25mOhm
L_X20Y100VDD_X20Y110VDD X20Y105VDD X20Y110VDD 2.91e-06nH
R_X20Y100VSS_X20Y110VSS X20Y100VSS X20Y105VSS 25mOhm
L_X20Y100VSS_X20Y110VSS X20Y105VSS X20Y110VSS 2.91e-06nH
R_X20Y110VDD_X20Y120VDD X20Y110VDD X20Y115VDD 25mOhm
L_X20Y110VDD_X20Y120VDD X20Y115VDD X20Y120VDD 2.91e-06nH
R_X20Y110VSS_X20Y120VSS X20Y110VSS X20Y115VSS 25mOhm
L_X20Y110VSS_X20Y120VSS X20Y115VSS X20Y120VSS 2.91e-06nH
R_X30Y10VDD_X30Y20VDD X30Y10VDD X30Y15VDD 25mOhm
L_X30Y10VDD_X30Y20VDD X30Y15VDD X30Y20VDD 2.91e-06nH
R_X30Y10VSS_X30Y20VSS X30Y10VSS X30Y15VSS 25mOhm
L_X30Y10VSS_X30Y20VSS X30Y15VSS X30Y20VSS 2.91e-06nH
R_X30Y20VDD_X30Y30VDD X30Y20VDD X30Y25VDD 25mOhm
L_X30Y20VDD_X30Y30VDD X30Y25VDD X30Y30VDD 2.91e-06nH
R_X30Y20VSS_X30Y30VSS X30Y20VSS X30Y25VSS 25mOhm
L_X30Y20VSS_X30Y30VSS X30Y25VSS X30Y30VSS 2.91e-06nH
R_X30Y30VDD_X30Y40VDD X30Y30VDD X30Y35VDD 25mOhm
L_X30Y30VDD_X30Y40VDD X30Y35VDD X30Y40VDD 2.91e-06nH
R_X30Y30VSS_X30Y40VSS X30Y30VSS X30Y35VSS 25mOhm
L_X30Y30VSS_X30Y40VSS X30Y35VSS X30Y40VSS 2.91e-06nH
R_X30Y40VDD_X30Y50VDD X30Y40VDD X30Y45VDD 25mOhm
L_X30Y40VDD_X30Y50VDD X30Y45VDD X30Y50VDD 2.91e-06nH
R_X30Y40VSS_X30Y50VSS X30Y40VSS X30Y45VSS 25mOhm
L_X30Y40VSS_X30Y50VSS X30Y45VSS X30Y50VSS 2.91e-06nH
R_X30Y50VDD_X30Y60VDD X30Y50VDD X30Y55VDD 25mOhm
L_X30Y50VDD_X30Y60VDD X30Y55VDD X30Y60VDD 2.91e-06nH
R_X30Y50VSS_X30Y60VSS X30Y50VSS X30Y55VSS 25mOhm
L_X30Y50VSS_X30Y60VSS X30Y55VSS X30Y60VSS 2.91e-06nH
R_X30Y60VDD_X30Y70VDD X30Y60VDD X30Y65VDD 25mOhm
L_X30Y60VDD_X30Y70VDD X30Y65VDD X30Y70VDD 2.91e-06nH
R_X30Y60VSS_X30Y70VSS X30Y60VSS X30Y65VSS 25mOhm
L_X30Y60VSS_X30Y70VSS X30Y65VSS X30Y70VSS 2.91e-06nH
R_X30Y70VDD_X30Y80VDD X30Y70VDD X30Y75VDD 25mOhm
L_X30Y70VDD_X30Y80VDD X30Y75VDD X30Y80VDD 2.91e-06nH
R_X30Y70VSS_X30Y80VSS X30Y70VSS X30Y75VSS 25mOhm
L_X30Y70VSS_X30Y80VSS X30Y75VSS X30Y80VSS 2.91e-06nH
R_X30Y80VDD_X30Y90VDD X30Y80VDD X30Y85VDD 25mOhm
L_X30Y80VDD_X30Y90VDD X30Y85VDD X30Y90VDD 2.91e-06nH
R_X30Y80VSS_X30Y90VSS X30Y80VSS X30Y85VSS 25mOhm
L_X30Y80VSS_X30Y90VSS X30Y85VSS X30Y90VSS 2.91e-06nH
R_X30Y90VDD_X30Y100VDD X30Y90VDD X30Y95VDD 25mOhm
L_X30Y90VDD_X30Y100VDD X30Y95VDD X30Y100VDD 2.91e-06nH
R_X30Y90VSS_X30Y100VSS X30Y90VSS X30Y95VSS 25mOhm
L_X30Y90VSS_X30Y100VSS X30Y95VSS X30Y100VSS 2.91e-06nH
R_X30Y100VDD_X30Y110VDD X30Y100VDD X30Y105VDD 25mOhm
L_X30Y100VDD_X30Y110VDD X30Y105VDD X30Y110VDD 2.91e-06nH
R_X30Y100VSS_X30Y110VSS X30Y100VSS X30Y105VSS 25mOhm
L_X30Y100VSS_X30Y110VSS X30Y105VSS X30Y110VSS 2.91e-06nH
R_X30Y110VDD_X30Y120VDD X30Y110VDD X30Y115VDD 25mOhm
L_X30Y110VDD_X30Y120VDD X30Y115VDD X30Y120VDD 2.91e-06nH
R_X30Y110VSS_X30Y120VSS X30Y110VSS X30Y115VSS 25mOhm
L_X30Y110VSS_X30Y120VSS X30Y115VSS X30Y120VSS 2.91e-06nH
R_X40Y10VDD_X40Y20VDD X40Y10VDD X40Y15VDD 25mOhm
L_X40Y10VDD_X40Y20VDD X40Y15VDD X40Y20VDD 2.91e-06nH
R_X40Y10VSS_X40Y20VSS X40Y10VSS X40Y15VSS 25mOhm
L_X40Y10VSS_X40Y20VSS X40Y15VSS X40Y20VSS 2.91e-06nH
R_X40Y20VDD_X40Y30VDD X40Y20VDD X40Y25VDD 25mOhm
L_X40Y20VDD_X40Y30VDD X40Y25VDD X40Y30VDD 2.91e-06nH
R_X40Y20VSS_X40Y30VSS X40Y20VSS X40Y25VSS 25mOhm
L_X40Y20VSS_X40Y30VSS X40Y25VSS X40Y30VSS 2.91e-06nH
R_X40Y30VDD_X40Y40VDD X40Y30VDD X40Y35VDD 25mOhm
L_X40Y30VDD_X40Y40VDD X40Y35VDD X40Y40VDD 2.91e-06nH
R_X40Y30VSS_X40Y40VSS X40Y30VSS X40Y35VSS 25mOhm
L_X40Y30VSS_X40Y40VSS X40Y35VSS X40Y40VSS 2.91e-06nH
R_X40Y40VDD_X40Y50VDD X40Y40VDD X40Y45VDD 25mOhm
L_X40Y40VDD_X40Y50VDD X40Y45VDD X40Y50VDD 2.91e-06nH
R_X40Y40VSS_X40Y50VSS X40Y40VSS X40Y45VSS 25mOhm
L_X40Y40VSS_X40Y50VSS X40Y45VSS X40Y50VSS 2.91e-06nH
R_X40Y50VDD_X40Y60VDD X40Y50VDD X40Y55VDD 25mOhm
L_X40Y50VDD_X40Y60VDD X40Y55VDD X40Y60VDD 2.91e-06nH
R_X40Y50VSS_X40Y60VSS X40Y50VSS X40Y55VSS 25mOhm
L_X40Y50VSS_X40Y60VSS X40Y55VSS X40Y60VSS 2.91e-06nH
R_X40Y60VDD_X40Y70VDD X40Y60VDD X40Y65VDD 25mOhm
L_X40Y60VDD_X40Y70VDD X40Y65VDD X40Y70VDD 2.91e-06nH
R_X40Y60VSS_X40Y70VSS X40Y60VSS X40Y65VSS 25mOhm
L_X40Y60VSS_X40Y70VSS X40Y65VSS X40Y70VSS 2.91e-06nH
R_X40Y70VDD_X40Y80VDD X40Y70VDD X40Y75VDD 25mOhm
L_X40Y70VDD_X40Y80VDD X40Y75VDD X40Y80VDD 2.91e-06nH
R_X40Y70VSS_X40Y80VSS X40Y70VSS X40Y75VSS 25mOhm
L_X40Y70VSS_X40Y80VSS X40Y75VSS X40Y80VSS 2.91e-06nH
R_X40Y80VDD_X40Y90VDD X40Y80VDD X40Y85VDD 25mOhm
L_X40Y80VDD_X40Y90VDD X40Y85VDD X40Y90VDD 2.91e-06nH
R_X40Y80VSS_X40Y90VSS X40Y80VSS X40Y85VSS 25mOhm
L_X40Y80VSS_X40Y90VSS X40Y85VSS X40Y90VSS 2.91e-06nH
R_X40Y90VDD_X40Y100VDD X40Y90VDD X40Y95VDD 25mOhm
L_X40Y90VDD_X40Y100VDD X40Y95VDD X40Y100VDD 2.91e-06nH
R_X40Y90VSS_X40Y100VSS X40Y90VSS X40Y95VSS 25mOhm
L_X40Y90VSS_X40Y100VSS X40Y95VSS X40Y100VSS 2.91e-06nH
R_X40Y100VDD_X40Y110VDD X40Y100VDD X40Y105VDD 25mOhm
L_X40Y100VDD_X40Y110VDD X40Y105VDD X40Y110VDD 2.91e-06nH
R_X40Y100VSS_X40Y110VSS X40Y100VSS X40Y105VSS 25mOhm
L_X40Y100VSS_X40Y110VSS X40Y105VSS X40Y110VSS 2.91e-06nH
R_X40Y110VDD_X40Y120VDD X40Y110VDD X40Y115VDD 25mOhm
L_X40Y110VDD_X40Y120VDD X40Y115VDD X40Y120VDD 2.91e-06nH
R_X40Y110VSS_X40Y120VSS X40Y110VSS X40Y115VSS 25mOhm
L_X40Y110VSS_X40Y120VSS X40Y115VSS X40Y120VSS 2.91e-06nH
R_X50Y10VDD_X50Y20VDD X50Y10VDD X50Y15VDD 25mOhm
L_X50Y10VDD_X50Y20VDD X50Y15VDD X50Y20VDD 2.91e-06nH
R_X50Y10VSS_X50Y20VSS X50Y10VSS X50Y15VSS 25mOhm
L_X50Y10VSS_X50Y20VSS X50Y15VSS X50Y20VSS 2.91e-06nH
R_X50Y20VDD_X50Y30VDD X50Y20VDD X50Y25VDD 25mOhm
L_X50Y20VDD_X50Y30VDD X50Y25VDD X50Y30VDD 2.91e-06nH
R_X50Y20VSS_X50Y30VSS X50Y20VSS X50Y25VSS 25mOhm
L_X50Y20VSS_X50Y30VSS X50Y25VSS X50Y30VSS 2.91e-06nH
R_X50Y30VDD_X50Y40VDD X50Y30VDD X50Y35VDD 25mOhm
L_X50Y30VDD_X50Y40VDD X50Y35VDD X50Y40VDD 2.91e-06nH
R_X50Y30VSS_X50Y40VSS X50Y30VSS X50Y35VSS 25mOhm
L_X50Y30VSS_X50Y40VSS X50Y35VSS X50Y40VSS 2.91e-06nH
R_X50Y40VDD_X50Y50VDD X50Y40VDD X50Y45VDD 25mOhm
L_X50Y40VDD_X50Y50VDD X50Y45VDD X50Y50VDD 2.91e-06nH
R_X50Y40VSS_X50Y50VSS X50Y40VSS X50Y45VSS 25mOhm
L_X50Y40VSS_X50Y50VSS X50Y45VSS X50Y50VSS 2.91e-06nH
R_X50Y50VDD_X50Y60VDD X50Y50VDD X50Y55VDD 25mOhm
L_X50Y50VDD_X50Y60VDD X50Y55VDD X50Y60VDD 2.91e-06nH
R_X50Y50VSS_X50Y60VSS X50Y50VSS X50Y55VSS 25mOhm
L_X50Y50VSS_X50Y60VSS X50Y55VSS X50Y60VSS 2.91e-06nH
R_X50Y60VDD_X50Y70VDD X50Y60VDD X50Y65VDD 25mOhm
L_X50Y60VDD_X50Y70VDD X50Y65VDD X50Y70VDD 2.91e-06nH
R_X50Y60VSS_X50Y70VSS X50Y60VSS X50Y65VSS 25mOhm
L_X50Y60VSS_X50Y70VSS X50Y65VSS X50Y70VSS 2.91e-06nH
R_X50Y70VDD_X50Y80VDD X50Y70VDD X50Y75VDD 25mOhm
L_X50Y70VDD_X50Y80VDD X50Y75VDD X50Y80VDD 2.91e-06nH
R_X50Y70VSS_X50Y80VSS X50Y70VSS X50Y75VSS 25mOhm
L_X50Y70VSS_X50Y80VSS X50Y75VSS X50Y80VSS 2.91e-06nH
R_X50Y80VDD_X50Y90VDD X50Y80VDD X50Y85VDD 25mOhm
L_X50Y80VDD_X50Y90VDD X50Y85VDD X50Y90VDD 2.91e-06nH
R_X50Y80VSS_X50Y90VSS X50Y80VSS X50Y85VSS 25mOhm
L_X50Y80VSS_X50Y90VSS X50Y85VSS X50Y90VSS 2.91e-06nH
R_X50Y90VDD_X50Y100VDD X50Y90VDD X50Y95VDD 25mOhm
L_X50Y90VDD_X50Y100VDD X50Y95VDD X50Y100VDD 2.91e-06nH
R_X50Y90VSS_X50Y100VSS X50Y90VSS X50Y95VSS 25mOhm
L_X50Y90VSS_X50Y100VSS X50Y95VSS X50Y100VSS 2.91e-06nH
R_X50Y100VDD_X50Y110VDD X50Y100VDD X50Y105VDD 25mOhm
L_X50Y100VDD_X50Y110VDD X50Y105VDD X50Y110VDD 2.91e-06nH
R_X50Y100VSS_X50Y110VSS X50Y100VSS X50Y105VSS 25mOhm
L_X50Y100VSS_X50Y110VSS X50Y105VSS X50Y110VSS 2.91e-06nH
R_X50Y110VDD_X50Y120VDD X50Y110VDD X50Y115VDD 25mOhm
L_X50Y110VDD_X50Y120VDD X50Y115VDD X50Y120VDD 2.91e-06nH
R_X50Y110VSS_X50Y120VSS X50Y110VSS X50Y115VSS 25mOhm
L_X50Y110VSS_X50Y120VSS X50Y115VSS X50Y120VSS 2.91e-06nH
R_X60Y10VDD_X60Y20VDD X60Y10VDD X60Y15VDD 25mOhm
L_X60Y10VDD_X60Y20VDD X60Y15VDD X60Y20VDD 2.91e-06nH
R_X60Y10VSS_X60Y20VSS X60Y10VSS X60Y15VSS 25mOhm
L_X60Y10VSS_X60Y20VSS X60Y15VSS X60Y20VSS 2.91e-06nH
R_X60Y20VDD_X60Y30VDD X60Y20VDD X60Y25VDD 25mOhm
L_X60Y20VDD_X60Y30VDD X60Y25VDD X60Y30VDD 2.91e-06nH
R_X60Y20VSS_X60Y30VSS X60Y20VSS X60Y25VSS 25mOhm
L_X60Y20VSS_X60Y30VSS X60Y25VSS X60Y30VSS 2.91e-06nH
R_X60Y30VDD_X60Y40VDD X60Y30VDD X60Y35VDD 25mOhm
L_X60Y30VDD_X60Y40VDD X60Y35VDD X60Y40VDD 2.91e-06nH
R_X60Y30VSS_X60Y40VSS X60Y30VSS X60Y35VSS 25mOhm
L_X60Y30VSS_X60Y40VSS X60Y35VSS X60Y40VSS 2.91e-06nH
R_X60Y40VDD_X60Y50VDD X60Y40VDD X60Y45VDD 25mOhm
L_X60Y40VDD_X60Y50VDD X60Y45VDD X60Y50VDD 2.91e-06nH
R_X60Y40VSS_X60Y50VSS X60Y40VSS X60Y45VSS 25mOhm
L_X60Y40VSS_X60Y50VSS X60Y45VSS X60Y50VSS 2.91e-06nH
R_X60Y50VDD_X60Y60VDD X60Y50VDD X60Y55VDD 25mOhm
L_X60Y50VDD_X60Y60VDD X60Y55VDD X60Y60VDD 2.91e-06nH
R_X60Y50VSS_X60Y60VSS X60Y50VSS X60Y55VSS 25mOhm
L_X60Y50VSS_X60Y60VSS X60Y55VSS X60Y60VSS 2.91e-06nH
R_X60Y60VDD_X60Y70VDD X60Y60VDD X60Y65VDD 25mOhm
L_X60Y60VDD_X60Y70VDD X60Y65VDD X60Y70VDD 2.91e-06nH
R_X60Y60VSS_X60Y70VSS X60Y60VSS X60Y65VSS 25mOhm
L_X60Y60VSS_X60Y70VSS X60Y65VSS X60Y70VSS 2.91e-06nH
R_X60Y70VDD_X60Y80VDD X60Y70VDD X60Y75VDD 25mOhm
L_X60Y70VDD_X60Y80VDD X60Y75VDD X60Y80VDD 2.91e-06nH
R_X60Y70VSS_X60Y80VSS X60Y70VSS X60Y75VSS 25mOhm
L_X60Y70VSS_X60Y80VSS X60Y75VSS X60Y80VSS 2.91e-06nH
R_X60Y80VDD_X60Y90VDD X60Y80VDD X60Y85VDD 25mOhm
L_X60Y80VDD_X60Y90VDD X60Y85VDD X60Y90VDD 2.91e-06nH
R_X60Y80VSS_X60Y90VSS X60Y80VSS X60Y85VSS 25mOhm
L_X60Y80VSS_X60Y90VSS X60Y85VSS X60Y90VSS 2.91e-06nH
R_X60Y90VDD_X60Y100VDD X60Y90VDD X60Y95VDD 25mOhm
L_X60Y90VDD_X60Y100VDD X60Y95VDD X60Y100VDD 2.91e-06nH
R_X60Y90VSS_X60Y100VSS X60Y90VSS X60Y95VSS 25mOhm
L_X60Y90VSS_X60Y100VSS X60Y95VSS X60Y100VSS 2.91e-06nH
R_X60Y100VDD_X60Y110VDD X60Y100VDD X60Y105VDD 25mOhm
L_X60Y100VDD_X60Y110VDD X60Y105VDD X60Y110VDD 2.91e-06nH
R_X60Y100VSS_X60Y110VSS X60Y100VSS X60Y105VSS 25mOhm
L_X60Y100VSS_X60Y110VSS X60Y105VSS X60Y110VSS 2.91e-06nH
R_X60Y110VDD_X60Y120VDD X60Y110VDD X60Y115VDD 25mOhm
L_X60Y110VDD_X60Y120VDD X60Y115VDD X60Y120VDD 2.91e-06nH
R_X60Y110VSS_X60Y120VSS X60Y110VSS X60Y115VSS 25mOhm
L_X60Y110VSS_X60Y120VSS X60Y115VSS X60Y120VSS 2.91e-06nH
R_X70Y10VDD_X70Y20VDD X70Y10VDD X70Y15VDD 25mOhm
L_X70Y10VDD_X70Y20VDD X70Y15VDD X70Y20VDD 2.91e-06nH
R_X70Y10VSS_X70Y20VSS X70Y10VSS X70Y15VSS 25mOhm
L_X70Y10VSS_X70Y20VSS X70Y15VSS X70Y20VSS 2.91e-06nH
R_X70Y20VDD_X70Y30VDD X70Y20VDD X70Y25VDD 25mOhm
L_X70Y20VDD_X70Y30VDD X70Y25VDD X70Y30VDD 2.91e-06nH
R_X70Y20VSS_X70Y30VSS X70Y20VSS X70Y25VSS 25mOhm
L_X70Y20VSS_X70Y30VSS X70Y25VSS X70Y30VSS 2.91e-06nH
R_X70Y30VDD_X70Y40VDD X70Y30VDD X70Y35VDD 25mOhm
L_X70Y30VDD_X70Y40VDD X70Y35VDD X70Y40VDD 2.91e-06nH
R_X70Y30VSS_X70Y40VSS X70Y30VSS X70Y35VSS 25mOhm
L_X70Y30VSS_X70Y40VSS X70Y35VSS X70Y40VSS 2.91e-06nH
R_X70Y40VDD_X70Y50VDD X70Y40VDD X70Y45VDD 25mOhm
L_X70Y40VDD_X70Y50VDD X70Y45VDD X70Y50VDD 2.91e-06nH
R_X70Y40VSS_X70Y50VSS X70Y40VSS X70Y45VSS 25mOhm
L_X70Y40VSS_X70Y50VSS X70Y45VSS X70Y50VSS 2.91e-06nH
R_X70Y50VDD_X70Y60VDD X70Y50VDD X70Y55VDD 25mOhm
L_X70Y50VDD_X70Y60VDD X70Y55VDD X70Y60VDD 2.91e-06nH
R_X70Y50VSS_X70Y60VSS X70Y50VSS X70Y55VSS 25mOhm
L_X70Y50VSS_X70Y60VSS X70Y55VSS X70Y60VSS 2.91e-06nH
R_X70Y60VDD_X70Y70VDD X70Y60VDD X70Y65VDD 25mOhm
L_X70Y60VDD_X70Y70VDD X70Y65VDD X70Y70VDD 2.91e-06nH
R_X70Y60VSS_X70Y70VSS X70Y60VSS X70Y65VSS 25mOhm
L_X70Y60VSS_X70Y70VSS X70Y65VSS X70Y70VSS 2.91e-06nH
R_X70Y70VDD_X70Y80VDD X70Y70VDD X70Y75VDD 25mOhm
L_X70Y70VDD_X70Y80VDD X70Y75VDD X70Y80VDD 2.91e-06nH
R_X70Y70VSS_X70Y80VSS X70Y70VSS X70Y75VSS 25mOhm
L_X70Y70VSS_X70Y80VSS X70Y75VSS X70Y80VSS 2.91e-06nH
R_X70Y80VDD_X70Y90VDD X70Y80VDD X70Y85VDD 25mOhm
L_X70Y80VDD_X70Y90VDD X70Y85VDD X70Y90VDD 2.91e-06nH
R_X70Y80VSS_X70Y90VSS X70Y80VSS X70Y85VSS 25mOhm
L_X70Y80VSS_X70Y90VSS X70Y85VSS X70Y90VSS 2.91e-06nH
R_X70Y90VDD_X70Y100VDD X70Y90VDD X70Y95VDD 25mOhm
L_X70Y90VDD_X70Y100VDD X70Y95VDD X70Y100VDD 2.91e-06nH
R_X70Y90VSS_X70Y100VSS X70Y90VSS X70Y95VSS 25mOhm
L_X70Y90VSS_X70Y100VSS X70Y95VSS X70Y100VSS 2.91e-06nH
R_X70Y100VDD_X70Y110VDD X70Y100VDD X70Y105VDD 25mOhm
L_X70Y100VDD_X70Y110VDD X70Y105VDD X70Y110VDD 2.91e-06nH
R_X70Y100VSS_X70Y110VSS X70Y100VSS X70Y105VSS 25mOhm
L_X70Y100VSS_X70Y110VSS X70Y105VSS X70Y110VSS 2.91e-06nH
R_X70Y110VDD_X70Y120VDD X70Y110VDD X70Y115VDD 25mOhm
L_X70Y110VDD_X70Y120VDD X70Y115VDD X70Y120VDD 2.91e-06nH
R_X70Y110VSS_X70Y120VSS X70Y110VSS X70Y115VSS 25mOhm
L_X70Y110VSS_X70Y120VSS X70Y115VSS X70Y120VSS 2.91e-06nH
R_X80Y10VDD_X80Y20VDD X80Y10VDD X80Y15VDD 25mOhm
L_X80Y10VDD_X80Y20VDD X80Y15VDD X80Y20VDD 2.91e-06nH
R_X80Y10VSS_X80Y20VSS X80Y10VSS X80Y15VSS 25mOhm
L_X80Y10VSS_X80Y20VSS X80Y15VSS X80Y20VSS 2.91e-06nH
R_X80Y20VDD_X80Y30VDD X80Y20VDD X80Y25VDD 25mOhm
L_X80Y20VDD_X80Y30VDD X80Y25VDD X80Y30VDD 2.91e-06nH
R_X80Y20VSS_X80Y30VSS X80Y20VSS X80Y25VSS 25mOhm
L_X80Y20VSS_X80Y30VSS X80Y25VSS X80Y30VSS 2.91e-06nH
R_X80Y30VDD_X80Y40VDD X80Y30VDD X80Y35VDD 25mOhm
L_X80Y30VDD_X80Y40VDD X80Y35VDD X80Y40VDD 2.91e-06nH
R_X80Y30VSS_X80Y40VSS X80Y30VSS X80Y35VSS 25mOhm
L_X80Y30VSS_X80Y40VSS X80Y35VSS X80Y40VSS 2.91e-06nH
R_X80Y40VDD_X80Y50VDD X80Y40VDD X80Y45VDD 25mOhm
L_X80Y40VDD_X80Y50VDD X80Y45VDD X80Y50VDD 2.91e-06nH
R_X80Y40VSS_X80Y50VSS X80Y40VSS X80Y45VSS 25mOhm
L_X80Y40VSS_X80Y50VSS X80Y45VSS X80Y50VSS 2.91e-06nH
R_X80Y50VDD_X80Y60VDD X80Y50VDD X80Y55VDD 25mOhm
L_X80Y50VDD_X80Y60VDD X80Y55VDD X80Y60VDD 2.91e-06nH
R_X80Y50VSS_X80Y60VSS X80Y50VSS X80Y55VSS 25mOhm
L_X80Y50VSS_X80Y60VSS X80Y55VSS X80Y60VSS 2.91e-06nH
R_X80Y60VDD_X80Y70VDD X80Y60VDD X80Y65VDD 25mOhm
L_X80Y60VDD_X80Y70VDD X80Y65VDD X80Y70VDD 2.91e-06nH
R_X80Y60VSS_X80Y70VSS X80Y60VSS X80Y65VSS 25mOhm
L_X80Y60VSS_X80Y70VSS X80Y65VSS X80Y70VSS 2.91e-06nH
R_X80Y70VDD_X80Y80VDD X80Y70VDD X80Y75VDD 25mOhm
L_X80Y70VDD_X80Y80VDD X80Y75VDD X80Y80VDD 2.91e-06nH
R_X80Y70VSS_X80Y80VSS X80Y70VSS X80Y75VSS 25mOhm
L_X80Y70VSS_X80Y80VSS X80Y75VSS X80Y80VSS 2.91e-06nH
R_X80Y80VDD_X80Y90VDD X80Y80VDD X80Y85VDD 25mOhm
L_X80Y80VDD_X80Y90VDD X80Y85VDD X80Y90VDD 2.91e-06nH
R_X80Y80VSS_X80Y90VSS X80Y80VSS X80Y85VSS 25mOhm
L_X80Y80VSS_X80Y90VSS X80Y85VSS X80Y90VSS 2.91e-06nH
R_X80Y90VDD_X80Y100VDD X80Y90VDD X80Y95VDD 25mOhm
L_X80Y90VDD_X80Y100VDD X80Y95VDD X80Y100VDD 2.91e-06nH
R_X80Y90VSS_X80Y100VSS X80Y90VSS X80Y95VSS 25mOhm
L_X80Y90VSS_X80Y100VSS X80Y95VSS X80Y100VSS 2.91e-06nH
R_X80Y100VDD_X80Y110VDD X80Y100VDD X80Y105VDD 25mOhm
L_X80Y100VDD_X80Y110VDD X80Y105VDD X80Y110VDD 2.91e-06nH
R_X80Y100VSS_X80Y110VSS X80Y100VSS X80Y105VSS 25mOhm
L_X80Y100VSS_X80Y110VSS X80Y105VSS X80Y110VSS 2.91e-06nH
R_X80Y110VDD_X80Y120VDD X80Y110VDD X80Y115VDD 25mOhm
L_X80Y110VDD_X80Y120VDD X80Y115VDD X80Y120VDD 2.91e-06nH
R_X80Y110VSS_X80Y120VSS X80Y110VSS X80Y115VSS 25mOhm
L_X80Y110VSS_X80Y120VSS X80Y115VSS X80Y120VSS 2.91e-06nH
R_X90Y10VDD_X90Y20VDD X90Y10VDD X90Y15VDD 25mOhm
L_X90Y10VDD_X90Y20VDD X90Y15VDD X90Y20VDD 2.91e-06nH
R_X90Y10VSS_X90Y20VSS X90Y10VSS X90Y15VSS 25mOhm
L_X90Y10VSS_X90Y20VSS X90Y15VSS X90Y20VSS 2.91e-06nH
R_X90Y20VDD_X90Y30VDD X90Y20VDD X90Y25VDD 25mOhm
L_X90Y20VDD_X90Y30VDD X90Y25VDD X90Y30VDD 2.91e-06nH
R_X90Y20VSS_X90Y30VSS X90Y20VSS X90Y25VSS 25mOhm
L_X90Y20VSS_X90Y30VSS X90Y25VSS X90Y30VSS 2.91e-06nH
R_X90Y30VDD_X90Y40VDD X90Y30VDD X90Y35VDD 25mOhm
L_X90Y30VDD_X90Y40VDD X90Y35VDD X90Y40VDD 2.91e-06nH
R_X90Y30VSS_X90Y40VSS X90Y30VSS X90Y35VSS 25mOhm
L_X90Y30VSS_X90Y40VSS X90Y35VSS X90Y40VSS 2.91e-06nH
R_X90Y40VDD_X90Y50VDD X90Y40VDD X90Y45VDD 25mOhm
L_X90Y40VDD_X90Y50VDD X90Y45VDD X90Y50VDD 2.91e-06nH
R_X90Y40VSS_X90Y50VSS X90Y40VSS X90Y45VSS 25mOhm
L_X90Y40VSS_X90Y50VSS X90Y45VSS X90Y50VSS 2.91e-06nH
R_X90Y50VDD_X90Y60VDD X90Y50VDD X90Y55VDD 25mOhm
L_X90Y50VDD_X90Y60VDD X90Y55VDD X90Y60VDD 2.91e-06nH
R_X90Y50VSS_X90Y60VSS X90Y50VSS X90Y55VSS 25mOhm
L_X90Y50VSS_X90Y60VSS X90Y55VSS X90Y60VSS 2.91e-06nH
R_X90Y60VDD_X90Y70VDD X90Y60VDD X90Y65VDD 25mOhm
L_X90Y60VDD_X90Y70VDD X90Y65VDD X90Y70VDD 2.91e-06nH
R_X90Y60VSS_X90Y70VSS X90Y60VSS X90Y65VSS 25mOhm
L_X90Y60VSS_X90Y70VSS X90Y65VSS X90Y70VSS 2.91e-06nH
R_X90Y70VDD_X90Y80VDD X90Y70VDD X90Y75VDD 25mOhm
L_X90Y70VDD_X90Y80VDD X90Y75VDD X90Y80VDD 2.91e-06nH
R_X90Y70VSS_X90Y80VSS X90Y70VSS X90Y75VSS 25mOhm
L_X90Y70VSS_X90Y80VSS X90Y75VSS X90Y80VSS 2.91e-06nH
R_X90Y80VDD_X90Y90VDD X90Y80VDD X90Y85VDD 25mOhm
L_X90Y80VDD_X90Y90VDD X90Y85VDD X90Y90VDD 2.91e-06nH
R_X90Y80VSS_X90Y90VSS X90Y80VSS X90Y85VSS 25mOhm
L_X90Y80VSS_X90Y90VSS X90Y85VSS X90Y90VSS 2.91e-06nH
R_X90Y90VDD_X90Y100VDD X90Y90VDD X90Y95VDD 25mOhm
L_X90Y90VDD_X90Y100VDD X90Y95VDD X90Y100VDD 2.91e-06nH
R_X90Y90VSS_X90Y100VSS X90Y90VSS X90Y95VSS 25mOhm
L_X90Y90VSS_X90Y100VSS X90Y95VSS X90Y100VSS 2.91e-06nH
R_X90Y100VDD_X90Y110VDD X90Y100VDD X90Y105VDD 25mOhm
L_X90Y100VDD_X90Y110VDD X90Y105VDD X90Y110VDD 2.91e-06nH
R_X90Y100VSS_X90Y110VSS X90Y100VSS X90Y105VSS 25mOhm
L_X90Y100VSS_X90Y110VSS X90Y105VSS X90Y110VSS 2.91e-06nH
R_X90Y110VDD_X90Y120VDD X90Y110VDD X90Y115VDD 25mOhm
L_X90Y110VDD_X90Y120VDD X90Y115VDD X90Y120VDD 2.91e-06nH
R_X90Y110VSS_X90Y120VSS X90Y110VSS X90Y115VSS 25mOhm
L_X90Y110VSS_X90Y120VSS X90Y115VSS X90Y120VSS 2.91e-06nH
R_X100Y10VDD_X100Y20VDD X100Y10VDD X100Y15VDD 25mOhm
L_X100Y10VDD_X100Y20VDD X100Y15VDD X100Y20VDD 2.91e-06nH
R_X100Y10VSS_X100Y20VSS X100Y10VSS X100Y15VSS 25mOhm
L_X100Y10VSS_X100Y20VSS X100Y15VSS X100Y20VSS 2.91e-06nH
R_X100Y20VDD_X100Y30VDD X100Y20VDD X100Y25VDD 25mOhm
L_X100Y20VDD_X100Y30VDD X100Y25VDD X100Y30VDD 2.91e-06nH
R_X100Y20VSS_X100Y30VSS X100Y20VSS X100Y25VSS 25mOhm
L_X100Y20VSS_X100Y30VSS X100Y25VSS X100Y30VSS 2.91e-06nH
R_X100Y30VDD_X100Y40VDD X100Y30VDD X100Y35VDD 25mOhm
L_X100Y30VDD_X100Y40VDD X100Y35VDD X100Y40VDD 2.91e-06nH
R_X100Y30VSS_X100Y40VSS X100Y30VSS X100Y35VSS 25mOhm
L_X100Y30VSS_X100Y40VSS X100Y35VSS X100Y40VSS 2.91e-06nH
R_X100Y40VDD_X100Y50VDD X100Y40VDD X100Y45VDD 25mOhm
L_X100Y40VDD_X100Y50VDD X100Y45VDD X100Y50VDD 2.91e-06nH
R_X100Y40VSS_X100Y50VSS X100Y40VSS X100Y45VSS 25mOhm
L_X100Y40VSS_X100Y50VSS X100Y45VSS X100Y50VSS 2.91e-06nH
R_X100Y50VDD_X100Y60VDD X100Y50VDD X100Y55VDD 25mOhm
L_X100Y50VDD_X100Y60VDD X100Y55VDD X100Y60VDD 2.91e-06nH
R_X100Y50VSS_X100Y60VSS X100Y50VSS X100Y55VSS 25mOhm
L_X100Y50VSS_X100Y60VSS X100Y55VSS X100Y60VSS 2.91e-06nH
R_X100Y60VDD_X100Y70VDD X100Y60VDD X100Y65VDD 25mOhm
L_X100Y60VDD_X100Y70VDD X100Y65VDD X100Y70VDD 2.91e-06nH
R_X100Y60VSS_X100Y70VSS X100Y60VSS X100Y65VSS 25mOhm
L_X100Y60VSS_X100Y70VSS X100Y65VSS X100Y70VSS 2.91e-06nH
R_X100Y70VDD_X100Y80VDD X100Y70VDD X100Y75VDD 25mOhm
L_X100Y70VDD_X100Y80VDD X100Y75VDD X100Y80VDD 2.91e-06nH
R_X100Y70VSS_X100Y80VSS X100Y70VSS X100Y75VSS 25mOhm
L_X100Y70VSS_X100Y80VSS X100Y75VSS X100Y80VSS 2.91e-06nH
R_X100Y80VDD_X100Y90VDD X100Y80VDD X100Y85VDD 25mOhm
L_X100Y80VDD_X100Y90VDD X100Y85VDD X100Y90VDD 2.91e-06nH
R_X100Y80VSS_X100Y90VSS X100Y80VSS X100Y85VSS 25mOhm
L_X100Y80VSS_X100Y90VSS X100Y85VSS X100Y90VSS 2.91e-06nH
R_X100Y90VDD_X100Y100VDD X100Y90VDD X100Y95VDD 25mOhm
L_X100Y90VDD_X100Y100VDD X100Y95VDD X100Y100VDD 2.91e-06nH
R_X100Y90VSS_X100Y100VSS X100Y90VSS X100Y95VSS 25mOhm
L_X100Y90VSS_X100Y100VSS X100Y95VSS X100Y100VSS 2.91e-06nH
R_X100Y100VDD_X100Y110VDD X100Y100VDD X100Y105VDD 25mOhm
L_X100Y100VDD_X100Y110VDD X100Y105VDD X100Y110VDD 2.91e-06nH
R_X100Y100VSS_X100Y110VSS X100Y100VSS X100Y105VSS 25mOhm
L_X100Y100VSS_X100Y110VSS X100Y105VSS X100Y110VSS 2.91e-06nH
R_X100Y110VDD_X100Y120VDD X100Y110VDD X100Y115VDD 25mOhm
L_X100Y110VDD_X100Y120VDD X100Y115VDD X100Y120VDD 2.91e-06nH
R_X100Y110VSS_X100Y120VSS X100Y110VSS X100Y115VSS 25mOhm
L_X100Y110VSS_X100Y120VSS X100Y115VSS X100Y120VSS 2.91e-06nH
R_X110Y10VDD_X110Y20VDD X110Y10VDD X110Y15VDD 25mOhm
L_X110Y10VDD_X110Y20VDD X110Y15VDD X110Y20VDD 2.91e-06nH
R_X110Y10VSS_X110Y20VSS X110Y10VSS X110Y15VSS 25mOhm
L_X110Y10VSS_X110Y20VSS X110Y15VSS X110Y20VSS 2.91e-06nH
R_X110Y20VDD_X110Y30VDD X110Y20VDD X110Y25VDD 25mOhm
L_X110Y20VDD_X110Y30VDD X110Y25VDD X110Y30VDD 2.91e-06nH
R_X110Y20VSS_X110Y30VSS X110Y20VSS X110Y25VSS 25mOhm
L_X110Y20VSS_X110Y30VSS X110Y25VSS X110Y30VSS 2.91e-06nH
R_X110Y30VDD_X110Y40VDD X110Y30VDD X110Y35VDD 25mOhm
L_X110Y30VDD_X110Y40VDD X110Y35VDD X110Y40VDD 2.91e-06nH
R_X110Y30VSS_X110Y40VSS X110Y30VSS X110Y35VSS 25mOhm
L_X110Y30VSS_X110Y40VSS X110Y35VSS X110Y40VSS 2.91e-06nH
R_X110Y40VDD_X110Y50VDD X110Y40VDD X110Y45VDD 25mOhm
L_X110Y40VDD_X110Y50VDD X110Y45VDD X110Y50VDD 2.91e-06nH
R_X110Y40VSS_X110Y50VSS X110Y40VSS X110Y45VSS 25mOhm
L_X110Y40VSS_X110Y50VSS X110Y45VSS X110Y50VSS 2.91e-06nH
R_X110Y50VDD_X110Y60VDD X110Y50VDD X110Y55VDD 25mOhm
L_X110Y50VDD_X110Y60VDD X110Y55VDD X110Y60VDD 2.91e-06nH
R_X110Y50VSS_X110Y60VSS X110Y50VSS X110Y55VSS 25mOhm
L_X110Y50VSS_X110Y60VSS X110Y55VSS X110Y60VSS 2.91e-06nH
R_X110Y60VDD_X110Y70VDD X110Y60VDD X110Y65VDD 25mOhm
L_X110Y60VDD_X110Y70VDD X110Y65VDD X110Y70VDD 2.91e-06nH
R_X110Y60VSS_X110Y70VSS X110Y60VSS X110Y65VSS 25mOhm
L_X110Y60VSS_X110Y70VSS X110Y65VSS X110Y70VSS 2.91e-06nH
R_X110Y70VDD_X110Y80VDD X110Y70VDD X110Y75VDD 25mOhm
L_X110Y70VDD_X110Y80VDD X110Y75VDD X110Y80VDD 2.91e-06nH
R_X110Y70VSS_X110Y80VSS X110Y70VSS X110Y75VSS 25mOhm
L_X110Y70VSS_X110Y80VSS X110Y75VSS X110Y80VSS 2.91e-06nH
R_X110Y80VDD_X110Y90VDD X110Y80VDD X110Y85VDD 25mOhm
L_X110Y80VDD_X110Y90VDD X110Y85VDD X110Y90VDD 2.91e-06nH
R_X110Y80VSS_X110Y90VSS X110Y80VSS X110Y85VSS 25mOhm
L_X110Y80VSS_X110Y90VSS X110Y85VSS X110Y90VSS 2.91e-06nH
R_X110Y90VDD_X110Y100VDD X110Y90VDD X110Y95VDD 25mOhm
L_X110Y90VDD_X110Y100VDD X110Y95VDD X110Y100VDD 2.91e-06nH
R_X110Y90VSS_X110Y100VSS X110Y90VSS X110Y95VSS 25mOhm
L_X110Y90VSS_X110Y100VSS X110Y95VSS X110Y100VSS 2.91e-06nH
R_X110Y100VDD_X110Y110VDD X110Y100VDD X110Y105VDD 25mOhm
L_X110Y100VDD_X110Y110VDD X110Y105VDD X110Y110VDD 2.91e-06nH
R_X110Y100VSS_X110Y110VSS X110Y100VSS X110Y105VSS 25mOhm
L_X110Y100VSS_X110Y110VSS X110Y105VSS X110Y110VSS 2.91e-06nH
R_X110Y110VDD_X110Y120VDD X110Y110VDD X110Y115VDD 25mOhm
L_X110Y110VDD_X110Y120VDD X110Y115VDD X110Y120VDD 2.91e-06nH
R_X110Y110VSS_X110Y120VSS X110Y110VSS X110Y115VSS 25mOhm
L_X110Y110VSS_X110Y120VSS X110Y115VSS X110Y120VSS 2.91e-06nH
R_X120Y10VDD_X120Y20VDD X120Y10VDD X120Y15VDD 25mOhm
L_X120Y10VDD_X120Y20VDD X120Y15VDD X120Y20VDD 2.91e-06nH
R_X120Y10VSS_X120Y20VSS X120Y10VSS X120Y15VSS 25mOhm
L_X120Y10VSS_X120Y20VSS X120Y15VSS X120Y20VSS 2.91e-06nH
R_X120Y20VDD_X120Y30VDD X120Y20VDD X120Y25VDD 25mOhm
L_X120Y20VDD_X120Y30VDD X120Y25VDD X120Y30VDD 2.91e-06nH
R_X120Y20VSS_X120Y30VSS X120Y20VSS X120Y25VSS 25mOhm
L_X120Y20VSS_X120Y30VSS X120Y25VSS X120Y30VSS 2.91e-06nH
R_X120Y30VDD_X120Y40VDD X120Y30VDD X120Y35VDD 25mOhm
L_X120Y30VDD_X120Y40VDD X120Y35VDD X120Y40VDD 2.91e-06nH
R_X120Y30VSS_X120Y40VSS X120Y30VSS X120Y35VSS 25mOhm
L_X120Y30VSS_X120Y40VSS X120Y35VSS X120Y40VSS 2.91e-06nH
R_X120Y40VDD_X120Y50VDD X120Y40VDD X120Y45VDD 25mOhm
L_X120Y40VDD_X120Y50VDD X120Y45VDD X120Y50VDD 2.91e-06nH
R_X120Y40VSS_X120Y50VSS X120Y40VSS X120Y45VSS 25mOhm
L_X120Y40VSS_X120Y50VSS X120Y45VSS X120Y50VSS 2.91e-06nH
R_X120Y50VDD_X120Y60VDD X120Y50VDD X120Y55VDD 25mOhm
L_X120Y50VDD_X120Y60VDD X120Y55VDD X120Y60VDD 2.91e-06nH
R_X120Y50VSS_X120Y60VSS X120Y50VSS X120Y55VSS 25mOhm
L_X120Y50VSS_X120Y60VSS X120Y55VSS X120Y60VSS 2.91e-06nH
R_X120Y60VDD_X120Y70VDD X120Y60VDD X120Y65VDD 25mOhm
L_X120Y60VDD_X120Y70VDD X120Y65VDD X120Y70VDD 2.91e-06nH
R_X120Y60VSS_X120Y70VSS X120Y60VSS X120Y65VSS 25mOhm
L_X120Y60VSS_X120Y70VSS X120Y65VSS X120Y70VSS 2.91e-06nH
R_X120Y70VDD_X120Y80VDD X120Y70VDD X120Y75VDD 25mOhm
L_X120Y70VDD_X120Y80VDD X120Y75VDD X120Y80VDD 2.91e-06nH
R_X120Y70VSS_X120Y80VSS X120Y70VSS X120Y75VSS 25mOhm
L_X120Y70VSS_X120Y80VSS X120Y75VSS X120Y80VSS 2.91e-06nH
R_X120Y80VDD_X120Y90VDD X120Y80VDD X120Y85VDD 25mOhm
L_X120Y80VDD_X120Y90VDD X120Y85VDD X120Y90VDD 2.91e-06nH
R_X120Y80VSS_X120Y90VSS X120Y80VSS X120Y85VSS 25mOhm
L_X120Y80VSS_X120Y90VSS X120Y85VSS X120Y90VSS 2.91e-06nH
R_X120Y90VDD_X120Y100VDD X120Y90VDD X120Y95VDD 25mOhm
L_X120Y90VDD_X120Y100VDD X120Y95VDD X120Y100VDD 2.91e-06nH
R_X120Y90VSS_X120Y100VSS X120Y90VSS X120Y95VSS 25mOhm
L_X120Y90VSS_X120Y100VSS X120Y95VSS X120Y100VSS 2.91e-06nH
R_X120Y100VDD_X120Y110VDD X120Y100VDD X120Y105VDD 25mOhm
L_X120Y100VDD_X120Y110VDD X120Y105VDD X120Y110VDD 2.91e-06nH
R_X120Y100VSS_X120Y110VSS X120Y100VSS X120Y105VSS 25mOhm
L_X120Y100VSS_X120Y110VSS X120Y105VSS X120Y110VSS 2.91e-06nH
R_X120Y110VDD_X120Y120VDD X120Y110VDD X120Y115VDD 25mOhm
L_X120Y110VDD_X120Y120VDD X120Y115VDD X120Y120VDD 2.91e-06nH
R_X120Y110VSS_X120Y120VSS X120Y110VSS X120Y115VSS 25mOhm
L_X120Y110VSS_X120Y120VSS X120Y115VSS X120Y120VSS 2.91e-06nH
C_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VSS 10nF
C_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VSS 10nF
C_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VSS 10nF
C_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VSS 10nF
C_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VSS 10nF
C_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VSS 10nF
C_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VSS 10nF
C_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VSS 10nF
C_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VSS 10nF
C_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VSS 10nF
C_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VSS 10nF
C_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VSS 10nF
C_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VSS 10nF
C_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VSS 10nF
C_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VSS 10nF
C_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VSS 10nF
C_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VSS 10nF
C_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VSS 10nF
C_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VSS 10nF
C_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VSS 10nF
C_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VSS 10nF
C_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VSS 10nF
C_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VSS 10nF
C_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VSS 10nF
C_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VSS 10nF
C_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VSS 10nF
C_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VSS 10nF
C_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VSS 10nF
C_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VSS 10nF
C_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VSS 10nF
C_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VSS 10nF
C_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VSS 10nF
C_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VSS 10nF
C_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VSS 10nF
C_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VSS 10nF
C_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VSS 10nF
C_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VSS 10nF
C_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VSS 10nF
C_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VSS 10nF
C_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VSS 10nF
C_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VSS 10nF
C_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VSS 10nF
C_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VSS 10nF
C_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VSS 10nF
C_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VSS 10nF
C_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VSS 10nF
C_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VSS 10nF
C_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VSS 10nF
C_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VSS 10nF
C_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VSS 10nF
C_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VSS 10nF
C_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VSS 10nF
C_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VSS 10nF
C_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VSS 10nF
C_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VSS 10nF
C_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VSS 10nF
C_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VSS 10nF
C_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VSS 10nF
C_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VSS 10nF
C_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VSS 10nF
C_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VSS 10nF
C_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VSS 10nF
C_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VSS 10nF
C_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VSS 10nF
C_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VSS 10nF
C_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VSS 10nF
C_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VSS 10nF
C_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VSS 10nF
C_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VSS 10nF
C_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VSS 10nF
C_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VSS 10nF
C_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VSS 10nF
C_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VSS 10nF
C_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VSS 10nF
C_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VSS 10nF
C_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VSS 10nF
C_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VSS 10nF
C_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VSS 10nF
C_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VSS 10nF
C_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VSS 10nF
C_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VSS 10nF
C_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VSS 10nF
C_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VSS 10nF
C_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VSS 10nF
C_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VSS 10nF
C_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VSS 10nF
C_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VSS 10nF
C_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VSS 10nF
C_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VSS 10nF
C_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VSS 10nF
C_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VSS 10nF
C_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VSS 10nF
C_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VSS 10nF
C_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VSS 10nF
C_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VSS 10nF
C_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VSS 10nF
C_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VSS 10nF
C_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VSS 10nF
C_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VSS 10nF
C_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VSS 10nF
C_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VSS 10nF
C_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VSS 10nF
C_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VSS 10nF
C_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VSS 10nF
C_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VSS 10nF
C_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VSS 10nF
C_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VSS 10nF
C_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VSS 10nF
C_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VSS 10nF
C_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VSS 10nF
C_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VSS 10nF
C_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VSS 10nF
C_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VSS 10nF
C_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VSS 10nF
C_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VSS 10nF
C_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VSS 10nF
C_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VSS 10nF
C_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VSS 10nF
C_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VSS 10nF
C_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VSS 10nF
C_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VSS 10nF
C_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VSS 10nF
C_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VSS 10nF
C_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VSS 10nF
C_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VSS 10nF
C_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VSS 10nF
C_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VSS 10nF
C_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VSS 10nF
C_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VSS 10nF
C_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VSS 10nF
C_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VSS 10nF
C_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VSS 10nF
C_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VSS 10nF
C_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VSS 10nF
C_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VSS 10nF
C_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VSS 10nF
C_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VSS 10nF
C_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VSS 10nF
C_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VSS 10nF
C_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VSS 10nF
C_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VSS 10nF
C_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VSS 10nF
C_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VSS 10nF
C_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VSS 10nF
I_X120Y120VDD_X120Y120VSS X120Y120VDD X120Y120VDDDM 1 AC=0.006944444444444444
V_X120Y120VDD_X120Y120VSS X120Y120VDDDM X120Y120VSS 0
I_X120Y10VDD_X120Y10VSS X120Y10VDD X120Y10VDDDM 1 AC=0.006944444444444444
V_X120Y10VDD_X120Y10VSS X120Y10VDDDM X120Y10VSS 0
I_X120Y20VDD_X120Y20VSS X120Y20VDD X120Y20VDDDM 1 AC=0.006944444444444444
V_X120Y20VDD_X120Y20VSS X120Y20VDDDM X120Y20VSS 0
I_X120Y30VDD_X120Y30VSS X120Y30VDD X120Y30VDDDM 1 AC=0.006944444444444444
V_X120Y30VDD_X120Y30VSS X120Y30VDDDM X120Y30VSS 0
I_X120Y40VDD_X120Y40VSS X120Y40VDD X120Y40VDDDM 1 AC=0.006944444444444444
V_X120Y40VDD_X120Y40VSS X120Y40VDDDM X120Y40VSS 0
I_X120Y50VDD_X120Y50VSS X120Y50VDD X120Y50VDDDM 1 AC=0.006944444444444444
V_X120Y50VDD_X120Y50VSS X120Y50VDDDM X120Y50VSS 0
I_X120Y60VDD_X120Y60VSS X120Y60VDD X120Y60VDDDM 1 AC=0.006944444444444444
V_X120Y60VDD_X120Y60VSS X120Y60VDDDM X120Y60VSS 0
I_X120Y70VDD_X120Y70VSS X120Y70VDD X120Y70VDDDM 1 AC=0.006944444444444444
V_X120Y70VDD_X120Y70VSS X120Y70VDDDM X120Y70VSS 0
I_X120Y80VDD_X120Y80VSS X120Y80VDD X120Y80VDDDM 1 AC=0.006944444444444444
V_X120Y80VDD_X120Y80VSS X120Y80VDDDM X120Y80VSS 0
I_X120Y90VDD_X120Y90VSS X120Y90VDD X120Y90VDDDM 1 AC=0.006944444444444444
V_X120Y90VDD_X120Y90VSS X120Y90VDDDM X120Y90VSS 0
I_X120Y100VDD_X120Y100VSS X120Y100VDD X120Y100VDDDM 1 AC=0.006944444444444444
V_X120Y100VDD_X120Y100VSS X120Y100VDDDM X120Y100VSS 0
I_X120Y110VDD_X120Y110VSS X120Y110VDD X120Y110VDDDM 1 AC=0.006944444444444444
V_X120Y110VDD_X120Y110VSS X120Y110VDDDM X120Y110VSS 0
I_X10Y120VDD_X10Y120VSS X10Y120VDD X10Y120VDDDM 1 AC=0.006944444444444444
V_X10Y120VDD_X10Y120VSS X10Y120VDDDM X10Y120VSS 0
I_X10Y10VDD_X10Y10VSS X10Y10VDD X10Y10VDDDM 1 AC=0.006944444444444444
V_X10Y10VDD_X10Y10VSS X10Y10VDDDM X10Y10VSS 0
I_X10Y20VDD_X10Y20VSS X10Y20VDD X10Y20VDDDM 1 AC=0.006944444444444444
V_X10Y20VDD_X10Y20VSS X10Y20VDDDM X10Y20VSS 0
I_X10Y30VDD_X10Y30VSS X10Y30VDD X10Y30VDDDM 1 AC=0.006944444444444444
V_X10Y30VDD_X10Y30VSS X10Y30VDDDM X10Y30VSS 0
I_X10Y40VDD_X10Y40VSS X10Y40VDD X10Y40VDDDM 1 AC=0.006944444444444444
V_X10Y40VDD_X10Y40VSS X10Y40VDDDM X10Y40VSS 0
I_X10Y50VDD_X10Y50VSS X10Y50VDD X10Y50VDDDM 1 AC=0.006944444444444444
V_X10Y50VDD_X10Y50VSS X10Y50VDDDM X10Y50VSS 0
I_X10Y60VDD_X10Y60VSS X10Y60VDD X10Y60VDDDM 1 AC=0.006944444444444444
V_X10Y60VDD_X10Y60VSS X10Y60VDDDM X10Y60VSS 0
I_X10Y70VDD_X10Y70VSS X10Y70VDD X10Y70VDDDM 1 AC=0.006944444444444444
V_X10Y70VDD_X10Y70VSS X10Y70VDDDM X10Y70VSS 0
I_X10Y80VDD_X10Y80VSS X10Y80VDD X10Y80VDDDM 1 AC=0.006944444444444444
V_X10Y80VDD_X10Y80VSS X10Y80VDDDM X10Y80VSS 0
I_X10Y90VDD_X10Y90VSS X10Y90VDD X10Y90VDDDM 1 AC=0.006944444444444444
V_X10Y90VDD_X10Y90VSS X10Y90VDDDM X10Y90VSS 0
I_X10Y100VDD_X10Y100VSS X10Y100VDD X10Y100VDDDM 1 AC=0.006944444444444444
V_X10Y100VDD_X10Y100VSS X10Y100VDDDM X10Y100VSS 0
I_X10Y110VDD_X10Y110VSS X10Y110VDD X10Y110VDDDM 1 AC=0.006944444444444444
V_X10Y110VDD_X10Y110VSS X10Y110VDDDM X10Y110VSS 0
I_X20Y120VDD_X20Y120VSS X20Y120VDD X20Y120VDDDM 1 AC=0.006944444444444444
V_X20Y120VDD_X20Y120VSS X20Y120VDDDM X20Y120VSS 0
I_X20Y10VDD_X20Y10VSS X20Y10VDD X20Y10VDDDM 1 AC=0.006944444444444444
V_X20Y10VDD_X20Y10VSS X20Y10VDDDM X20Y10VSS 0
I_X20Y20VDD_X20Y20VSS X20Y20VDD X20Y20VDDDM 1 AC=0.006944444444444444
V_X20Y20VDD_X20Y20VSS X20Y20VDDDM X20Y20VSS 0
I_X20Y30VDD_X20Y30VSS X20Y30VDD X20Y30VDDDM 1 AC=0.006944444444444444
V_X20Y30VDD_X20Y30VSS X20Y30VDDDM X20Y30VSS 0
I_X20Y40VDD_X20Y40VSS X20Y40VDD X20Y40VDDDM 1 AC=0.006944444444444444
V_X20Y40VDD_X20Y40VSS X20Y40VDDDM X20Y40VSS 0
I_X20Y50VDD_X20Y50VSS X20Y50VDD X20Y50VDDDM 1 AC=0.006944444444444444
V_X20Y50VDD_X20Y50VSS X20Y50VDDDM X20Y50VSS 0
I_X20Y60VDD_X20Y60VSS X20Y60VDD X20Y60VDDDM 1 AC=0.006944444444444444
V_X20Y60VDD_X20Y60VSS X20Y60VDDDM X20Y60VSS 0
I_X20Y70VDD_X20Y70VSS X20Y70VDD X20Y70VDDDM 1 AC=0.006944444444444444
V_X20Y70VDD_X20Y70VSS X20Y70VDDDM X20Y70VSS 0
I_X20Y80VDD_X20Y80VSS X20Y80VDD X20Y80VDDDM 1 AC=0.006944444444444444
V_X20Y80VDD_X20Y80VSS X20Y80VDDDM X20Y80VSS 0
I_X20Y90VDD_X20Y90VSS X20Y90VDD X20Y90VDDDM 1 AC=0.006944444444444444
V_X20Y90VDD_X20Y90VSS X20Y90VDDDM X20Y90VSS 0
I_X20Y100VDD_X20Y100VSS X20Y100VDD X20Y100VDDDM 1 AC=0.006944444444444444
V_X20Y100VDD_X20Y100VSS X20Y100VDDDM X20Y100VSS 0
I_X20Y110VDD_X20Y110VSS X20Y110VDD X20Y110VDDDM 1 AC=0.006944444444444444
V_X20Y110VDD_X20Y110VSS X20Y110VDDDM X20Y110VSS 0
I_X30Y120VDD_X30Y120VSS X30Y120VDD X30Y120VDDDM 1 AC=0.006944444444444444
V_X30Y120VDD_X30Y120VSS X30Y120VDDDM X30Y120VSS 0
I_X30Y10VDD_X30Y10VSS X30Y10VDD X30Y10VDDDM 1 AC=0.006944444444444444
V_X30Y10VDD_X30Y10VSS X30Y10VDDDM X30Y10VSS 0
I_X30Y20VDD_X30Y20VSS X30Y20VDD X30Y20VDDDM 1 AC=0.006944444444444444
V_X30Y20VDD_X30Y20VSS X30Y20VDDDM X30Y20VSS 0
I_X30Y30VDD_X30Y30VSS X30Y30VDD X30Y30VDDDM 1 AC=0.006944444444444444
V_X30Y30VDD_X30Y30VSS X30Y30VDDDM X30Y30VSS 0
I_X30Y40VDD_X30Y40VSS X30Y40VDD X30Y40VDDDM 1 AC=0.006944444444444444
V_X30Y40VDD_X30Y40VSS X30Y40VDDDM X30Y40VSS 0
I_X30Y50VDD_X30Y50VSS X30Y50VDD X30Y50VDDDM 1 AC=0.006944444444444444
V_X30Y50VDD_X30Y50VSS X30Y50VDDDM X30Y50VSS 0
I_X30Y60VDD_X30Y60VSS X30Y60VDD X30Y60VDDDM 1 AC=0.006944444444444444
V_X30Y60VDD_X30Y60VSS X30Y60VDDDM X30Y60VSS 0
I_X30Y70VDD_X30Y70VSS X30Y70VDD X30Y70VDDDM 1 AC=0.006944444444444444
V_X30Y70VDD_X30Y70VSS X30Y70VDDDM X30Y70VSS 0
I_X30Y80VDD_X30Y80VSS X30Y80VDD X30Y80VDDDM 1 AC=0.006944444444444444
V_X30Y80VDD_X30Y80VSS X30Y80VDDDM X30Y80VSS 0
I_X30Y90VDD_X30Y90VSS X30Y90VDD X30Y90VDDDM 1 AC=0.006944444444444444
V_X30Y90VDD_X30Y90VSS X30Y90VDDDM X30Y90VSS 0
I_X30Y100VDD_X30Y100VSS X30Y100VDD X30Y100VDDDM 1 AC=0.006944444444444444
V_X30Y100VDD_X30Y100VSS X30Y100VDDDM X30Y100VSS 0
I_X30Y110VDD_X30Y110VSS X30Y110VDD X30Y110VDDDM 1 AC=0.006944444444444444
V_X30Y110VDD_X30Y110VSS X30Y110VDDDM X30Y110VSS 0
I_X40Y120VDD_X40Y120VSS X40Y120VDD X40Y120VDDDM 1 AC=0.006944444444444444
V_X40Y120VDD_X40Y120VSS X40Y120VDDDM X40Y120VSS 0
I_X40Y10VDD_X40Y10VSS X40Y10VDD X40Y10VDDDM 1 AC=0.006944444444444444
V_X40Y10VDD_X40Y10VSS X40Y10VDDDM X40Y10VSS 0
I_X40Y20VDD_X40Y20VSS X40Y20VDD X40Y20VDDDM 1 AC=0.006944444444444444
V_X40Y20VDD_X40Y20VSS X40Y20VDDDM X40Y20VSS 0
I_X40Y30VDD_X40Y30VSS X40Y30VDD X40Y30VDDDM 1 AC=0.006944444444444444
V_X40Y30VDD_X40Y30VSS X40Y30VDDDM X40Y30VSS 0
I_X40Y40VDD_X40Y40VSS X40Y40VDD X40Y40VDDDM 1 AC=0.006944444444444444
V_X40Y40VDD_X40Y40VSS X40Y40VDDDM X40Y40VSS 0
I_X40Y50VDD_X40Y50VSS X40Y50VDD X40Y50VDDDM 1 AC=0.006944444444444444
V_X40Y50VDD_X40Y50VSS X40Y50VDDDM X40Y50VSS 0
I_X40Y60VDD_X40Y60VSS X40Y60VDD X40Y60VDDDM 1 AC=0.006944444444444444
V_X40Y60VDD_X40Y60VSS X40Y60VDDDM X40Y60VSS 0
I_X40Y70VDD_X40Y70VSS X40Y70VDD X40Y70VDDDM 1 AC=0.006944444444444444
V_X40Y70VDD_X40Y70VSS X40Y70VDDDM X40Y70VSS 0
I_X40Y80VDD_X40Y80VSS X40Y80VDD X40Y80VDDDM 1 AC=0.006944444444444444
V_X40Y80VDD_X40Y80VSS X40Y80VDDDM X40Y80VSS 0
I_X40Y90VDD_X40Y90VSS X40Y90VDD X40Y90VDDDM 1 AC=0.006944444444444444
V_X40Y90VDD_X40Y90VSS X40Y90VDDDM X40Y90VSS 0
I_X40Y100VDD_X40Y100VSS X40Y100VDD X40Y100VDDDM 1 AC=0.006944444444444444
V_X40Y100VDD_X40Y100VSS X40Y100VDDDM X40Y100VSS 0
I_X40Y110VDD_X40Y110VSS X40Y110VDD X40Y110VDDDM 1 AC=0.006944444444444444
V_X40Y110VDD_X40Y110VSS X40Y110VDDDM X40Y110VSS 0
I_X50Y120VDD_X50Y120VSS X50Y120VDD X50Y120VDDDM 1 AC=0.006944444444444444
V_X50Y120VDD_X50Y120VSS X50Y120VDDDM X50Y120VSS 0
I_X50Y10VDD_X50Y10VSS X50Y10VDD X50Y10VDDDM 1 AC=0.006944444444444444
V_X50Y10VDD_X50Y10VSS X50Y10VDDDM X50Y10VSS 0
I_X50Y20VDD_X50Y20VSS X50Y20VDD X50Y20VDDDM 1 AC=0.006944444444444444
V_X50Y20VDD_X50Y20VSS X50Y20VDDDM X50Y20VSS 0
I_X50Y30VDD_X50Y30VSS X50Y30VDD X50Y30VDDDM 1 AC=0.006944444444444444
V_X50Y30VDD_X50Y30VSS X50Y30VDDDM X50Y30VSS 0
I_X50Y40VDD_X50Y40VSS X50Y40VDD X50Y40VDDDM 1 AC=0.006944444444444444
V_X50Y40VDD_X50Y40VSS X50Y40VDDDM X50Y40VSS 0
I_X50Y50VDD_X50Y50VSS X50Y50VDD X50Y50VDDDM 1 AC=0.006944444444444444
V_X50Y50VDD_X50Y50VSS X50Y50VDDDM X50Y50VSS 0
I_X50Y60VDD_X50Y60VSS X50Y60VDD X50Y60VDDDM 1 AC=0.006944444444444444
V_X50Y60VDD_X50Y60VSS X50Y60VDDDM X50Y60VSS 0
I_X50Y70VDD_X50Y70VSS X50Y70VDD X50Y70VDDDM 1 AC=0.006944444444444444
V_X50Y70VDD_X50Y70VSS X50Y70VDDDM X50Y70VSS 0
I_X50Y80VDD_X50Y80VSS X50Y80VDD X50Y80VDDDM 1 AC=0.006944444444444444
V_X50Y80VDD_X50Y80VSS X50Y80VDDDM X50Y80VSS 0
I_X50Y90VDD_X50Y90VSS X50Y90VDD X50Y90VDDDM 1 AC=0.006944444444444444
V_X50Y90VDD_X50Y90VSS X50Y90VDDDM X50Y90VSS 0
I_X50Y100VDD_X50Y100VSS X50Y100VDD X50Y100VDDDM 1 AC=0.006944444444444444
V_X50Y100VDD_X50Y100VSS X50Y100VDDDM X50Y100VSS 0
I_X50Y110VDD_X50Y110VSS X50Y110VDD X50Y110VDDDM 1 AC=0.006944444444444444
V_X50Y110VDD_X50Y110VSS X50Y110VDDDM X50Y110VSS 0
I_X60Y120VDD_X60Y120VSS X60Y120VDD X60Y120VDDDM 1 AC=0.006944444444444444
V_X60Y120VDD_X60Y120VSS X60Y120VDDDM X60Y120VSS 0
I_X60Y10VDD_X60Y10VSS X60Y10VDD X60Y10VDDDM 1 AC=0.006944444444444444
V_X60Y10VDD_X60Y10VSS X60Y10VDDDM X60Y10VSS 0
I_X60Y20VDD_X60Y20VSS X60Y20VDD X60Y20VDDDM 1 AC=0.006944444444444444
V_X60Y20VDD_X60Y20VSS X60Y20VDDDM X60Y20VSS 0
I_X60Y30VDD_X60Y30VSS X60Y30VDD X60Y30VDDDM 1 AC=0.006944444444444444
V_X60Y30VDD_X60Y30VSS X60Y30VDDDM X60Y30VSS 0
I_X60Y40VDD_X60Y40VSS X60Y40VDD X60Y40VDDDM 1 AC=0.006944444444444444
V_X60Y40VDD_X60Y40VSS X60Y40VDDDM X60Y40VSS 0
I_X60Y50VDD_X60Y50VSS X60Y50VDD X60Y50VDDDM 1 AC=0.006944444444444444
V_X60Y50VDD_X60Y50VSS X60Y50VDDDM X60Y50VSS 0
I_X60Y60VDD_X60Y60VSS X60Y60VDD X60Y60VDDDM 1 AC=0.006944444444444444
V_X60Y60VDD_X60Y60VSS X60Y60VDDDM X60Y60VSS 0
I_X60Y70VDD_X60Y70VSS X60Y70VDD X60Y70VDDDM 1 AC=0.006944444444444444
V_X60Y70VDD_X60Y70VSS X60Y70VDDDM X60Y70VSS 0
I_X60Y80VDD_X60Y80VSS X60Y80VDD X60Y80VDDDM 1 AC=0.006944444444444444
V_X60Y80VDD_X60Y80VSS X60Y80VDDDM X60Y80VSS 0
I_X60Y90VDD_X60Y90VSS X60Y90VDD X60Y90VDDDM 1 AC=0.006944444444444444
V_X60Y90VDD_X60Y90VSS X60Y90VDDDM X60Y90VSS 0
I_X60Y100VDD_X60Y100VSS X60Y100VDD X60Y100VDDDM 1 AC=0.006944444444444444
V_X60Y100VDD_X60Y100VSS X60Y100VDDDM X60Y100VSS 0
I_X60Y110VDD_X60Y110VSS X60Y110VDD X60Y110VDDDM 1 AC=0.006944444444444444
V_X60Y110VDD_X60Y110VSS X60Y110VDDDM X60Y110VSS 0
I_X70Y120VDD_X70Y120VSS X70Y120VDD X70Y120VDDDM 1 AC=0.006944444444444444
V_X70Y120VDD_X70Y120VSS X70Y120VDDDM X70Y120VSS 0
I_X70Y10VDD_X70Y10VSS X70Y10VDD X70Y10VDDDM 1 AC=0.006944444444444444
V_X70Y10VDD_X70Y10VSS X70Y10VDDDM X70Y10VSS 0
I_X70Y20VDD_X70Y20VSS X70Y20VDD X70Y20VDDDM 1 AC=0.006944444444444444
V_X70Y20VDD_X70Y20VSS X70Y20VDDDM X70Y20VSS 0
I_X70Y30VDD_X70Y30VSS X70Y30VDD X70Y30VDDDM 1 AC=0.006944444444444444
V_X70Y30VDD_X70Y30VSS X70Y30VDDDM X70Y30VSS 0
I_X70Y40VDD_X70Y40VSS X70Y40VDD X70Y40VDDDM 1 AC=0.006944444444444444
V_X70Y40VDD_X70Y40VSS X70Y40VDDDM X70Y40VSS 0
I_X70Y50VDD_X70Y50VSS X70Y50VDD X70Y50VDDDM 1 AC=0.006944444444444444
V_X70Y50VDD_X70Y50VSS X70Y50VDDDM X70Y50VSS 0
I_X70Y60VDD_X70Y60VSS X70Y60VDD X70Y60VDDDM 1 AC=0.006944444444444444
V_X70Y60VDD_X70Y60VSS X70Y60VDDDM X70Y60VSS 0
I_X70Y70VDD_X70Y70VSS X70Y70VDD X70Y70VDDDM 1 AC=0.006944444444444444
V_X70Y70VDD_X70Y70VSS X70Y70VDDDM X70Y70VSS 0
I_X70Y80VDD_X70Y80VSS X70Y80VDD X70Y80VDDDM 1 AC=0.006944444444444444
V_X70Y80VDD_X70Y80VSS X70Y80VDDDM X70Y80VSS 0
I_X70Y90VDD_X70Y90VSS X70Y90VDD X70Y90VDDDM 1 AC=0.006944444444444444
V_X70Y90VDD_X70Y90VSS X70Y90VDDDM X70Y90VSS 0
I_X70Y100VDD_X70Y100VSS X70Y100VDD X70Y100VDDDM 1 AC=0.006944444444444444
V_X70Y100VDD_X70Y100VSS X70Y100VDDDM X70Y100VSS 0
I_X70Y110VDD_X70Y110VSS X70Y110VDD X70Y110VDDDM 1 AC=0.006944444444444444
V_X70Y110VDD_X70Y110VSS X70Y110VDDDM X70Y110VSS 0
I_X80Y120VDD_X80Y120VSS X80Y120VDD X80Y120VDDDM 1 AC=0.006944444444444444
V_X80Y120VDD_X80Y120VSS X80Y120VDDDM X80Y120VSS 0
I_X80Y10VDD_X80Y10VSS X80Y10VDD X80Y10VDDDM 1 AC=0.006944444444444444
V_X80Y10VDD_X80Y10VSS X80Y10VDDDM X80Y10VSS 0
I_X80Y20VDD_X80Y20VSS X80Y20VDD X80Y20VDDDM 1 AC=0.006944444444444444
V_X80Y20VDD_X80Y20VSS X80Y20VDDDM X80Y20VSS 0
I_X80Y30VDD_X80Y30VSS X80Y30VDD X80Y30VDDDM 1 AC=0.006944444444444444
V_X80Y30VDD_X80Y30VSS X80Y30VDDDM X80Y30VSS 0
I_X80Y40VDD_X80Y40VSS X80Y40VDD X80Y40VDDDM 1 AC=0.006944444444444444
V_X80Y40VDD_X80Y40VSS X80Y40VDDDM X80Y40VSS 0
I_X80Y50VDD_X80Y50VSS X80Y50VDD X80Y50VDDDM 1 AC=0.006944444444444444
V_X80Y50VDD_X80Y50VSS X80Y50VDDDM X80Y50VSS 0
I_X80Y60VDD_X80Y60VSS X80Y60VDD X80Y60VDDDM 1 AC=0.006944444444444444
V_X80Y60VDD_X80Y60VSS X80Y60VDDDM X80Y60VSS 0
I_X80Y70VDD_X80Y70VSS X80Y70VDD X80Y70VDDDM 1 AC=0.006944444444444444
V_X80Y70VDD_X80Y70VSS X80Y70VDDDM X80Y70VSS 0
I_X80Y80VDD_X80Y80VSS X80Y80VDD X80Y80VDDDM 1 AC=0.006944444444444444
V_X80Y80VDD_X80Y80VSS X80Y80VDDDM X80Y80VSS 0
I_X80Y90VDD_X80Y90VSS X80Y90VDD X80Y90VDDDM 1 AC=0.006944444444444444
V_X80Y90VDD_X80Y90VSS X80Y90VDDDM X80Y90VSS 0
I_X80Y100VDD_X80Y100VSS X80Y100VDD X80Y100VDDDM 1 AC=0.006944444444444444
V_X80Y100VDD_X80Y100VSS X80Y100VDDDM X80Y100VSS 0
I_X80Y110VDD_X80Y110VSS X80Y110VDD X80Y110VDDDM 1 AC=0.006944444444444444
V_X80Y110VDD_X80Y110VSS X80Y110VDDDM X80Y110VSS 0
I_X90Y120VDD_X90Y120VSS X90Y120VDD X90Y120VDDDM 1 AC=0.006944444444444444
V_X90Y120VDD_X90Y120VSS X90Y120VDDDM X90Y120VSS 0
I_X90Y10VDD_X90Y10VSS X90Y10VDD X90Y10VDDDM 1 AC=0.006944444444444444
V_X90Y10VDD_X90Y10VSS X90Y10VDDDM X90Y10VSS 0
I_X90Y20VDD_X90Y20VSS X90Y20VDD X90Y20VDDDM 1 AC=0.006944444444444444
V_X90Y20VDD_X90Y20VSS X90Y20VDDDM X90Y20VSS 0
I_X90Y30VDD_X90Y30VSS X90Y30VDD X90Y30VDDDM 1 AC=0.006944444444444444
V_X90Y30VDD_X90Y30VSS X90Y30VDDDM X90Y30VSS 0
I_X90Y40VDD_X90Y40VSS X90Y40VDD X90Y40VDDDM 1 AC=0.006944444444444444
V_X90Y40VDD_X90Y40VSS X90Y40VDDDM X90Y40VSS 0
I_X90Y50VDD_X90Y50VSS X90Y50VDD X90Y50VDDDM 1 AC=0.006944444444444444
V_X90Y50VDD_X90Y50VSS X90Y50VDDDM X90Y50VSS 0
I_X90Y60VDD_X90Y60VSS X90Y60VDD X90Y60VDDDM 1 AC=0.006944444444444444
V_X90Y60VDD_X90Y60VSS X90Y60VDDDM X90Y60VSS 0
I_X90Y70VDD_X90Y70VSS X90Y70VDD X90Y70VDDDM 1 AC=0.006944444444444444
V_X90Y70VDD_X90Y70VSS X90Y70VDDDM X90Y70VSS 0
I_X90Y80VDD_X90Y80VSS X90Y80VDD X90Y80VDDDM 1 AC=0.006944444444444444
V_X90Y80VDD_X90Y80VSS X90Y80VDDDM X90Y80VSS 0
I_X90Y90VDD_X90Y90VSS X90Y90VDD X90Y90VDDDM 1 AC=0.006944444444444444
V_X90Y90VDD_X90Y90VSS X90Y90VDDDM X90Y90VSS 0
I_X90Y100VDD_X90Y100VSS X90Y100VDD X90Y100VDDDM 1 AC=0.006944444444444444
V_X90Y100VDD_X90Y100VSS X90Y100VDDDM X90Y100VSS 0
I_X90Y110VDD_X90Y110VSS X90Y110VDD X90Y110VDDDM 1 AC=0.006944444444444444
V_X90Y110VDD_X90Y110VSS X90Y110VDDDM X90Y110VSS 0
I_X100Y120VDD_X100Y120VSS X100Y120VDD X100Y120VDDDM 1 AC=0.006944444444444444
V_X100Y120VDD_X100Y120VSS X100Y120VDDDM X100Y120VSS 0
I_X100Y10VDD_X100Y10VSS X100Y10VDD X100Y10VDDDM 1 AC=0.006944444444444444
V_X100Y10VDD_X100Y10VSS X100Y10VDDDM X100Y10VSS 0
I_X100Y20VDD_X100Y20VSS X100Y20VDD X100Y20VDDDM 1 AC=0.006944444444444444
V_X100Y20VDD_X100Y20VSS X100Y20VDDDM X100Y20VSS 0
I_X100Y30VDD_X100Y30VSS X100Y30VDD X100Y30VDDDM 1 AC=0.006944444444444444
V_X100Y30VDD_X100Y30VSS X100Y30VDDDM X100Y30VSS 0
I_X100Y40VDD_X100Y40VSS X100Y40VDD X100Y40VDDDM 1 AC=0.006944444444444444
V_X100Y40VDD_X100Y40VSS X100Y40VDDDM X100Y40VSS 0
I_X100Y50VDD_X100Y50VSS X100Y50VDD X100Y50VDDDM 1 AC=0.006944444444444444
V_X100Y50VDD_X100Y50VSS X100Y50VDDDM X100Y50VSS 0
I_X100Y60VDD_X100Y60VSS X100Y60VDD X100Y60VDDDM 1 AC=0.006944444444444444
V_X100Y60VDD_X100Y60VSS X100Y60VDDDM X100Y60VSS 0
I_X100Y70VDD_X100Y70VSS X100Y70VDD X100Y70VDDDM 1 AC=0.006944444444444444
V_X100Y70VDD_X100Y70VSS X100Y70VDDDM X100Y70VSS 0
I_X100Y80VDD_X100Y80VSS X100Y80VDD X100Y80VDDDM 1 AC=0.006944444444444444
V_X100Y80VDD_X100Y80VSS X100Y80VDDDM X100Y80VSS 0
I_X100Y90VDD_X100Y90VSS X100Y90VDD X100Y90VDDDM 1 AC=0.006944444444444444
V_X100Y90VDD_X100Y90VSS X100Y90VDDDM X100Y90VSS 0
I_X100Y100VDD_X100Y100VSS X100Y100VDD X100Y100VDDDM 1 AC=0.006944444444444444
V_X100Y100VDD_X100Y100VSS X100Y100VDDDM X100Y100VSS 0
I_X100Y110VDD_X100Y110VSS X100Y110VDD X100Y110VDDDM 1 AC=0.006944444444444444
V_X100Y110VDD_X100Y110VSS X100Y110VDDDM X100Y110VSS 0
I_X110Y120VDD_X110Y120VSS X110Y120VDD X110Y120VDDDM 1 AC=0.006944444444444444
V_X110Y120VDD_X110Y120VSS X110Y120VDDDM X110Y120VSS 0
I_X110Y10VDD_X110Y10VSS X110Y10VDD X110Y10VDDDM 1 AC=0.006944444444444444
V_X110Y10VDD_X110Y10VSS X110Y10VDDDM X110Y10VSS 0
I_X110Y20VDD_X110Y20VSS X110Y20VDD X110Y20VDDDM 1 AC=0.006944444444444444
V_X110Y20VDD_X110Y20VSS X110Y20VDDDM X110Y20VSS 0
I_X110Y30VDD_X110Y30VSS X110Y30VDD X110Y30VDDDM 1 AC=0.006944444444444444
V_X110Y30VDD_X110Y30VSS X110Y30VDDDM X110Y30VSS 0
I_X110Y40VDD_X110Y40VSS X110Y40VDD X110Y40VDDDM 1 AC=0.006944444444444444
V_X110Y40VDD_X110Y40VSS X110Y40VDDDM X110Y40VSS 0
I_X110Y50VDD_X110Y50VSS X110Y50VDD X110Y50VDDDM 1 AC=0.006944444444444444
V_X110Y50VDD_X110Y50VSS X110Y50VDDDM X110Y50VSS 0
I_X110Y60VDD_X110Y60VSS X110Y60VDD X110Y60VDDDM 1 AC=0.006944444444444444
V_X110Y60VDD_X110Y60VSS X110Y60VDDDM X110Y60VSS 0
I_X110Y70VDD_X110Y70VSS X110Y70VDD X110Y70VDDDM 1 AC=0.006944444444444444
V_X110Y70VDD_X110Y70VSS X110Y70VDDDM X110Y70VSS 0
I_X110Y80VDD_X110Y80VSS X110Y80VDD X110Y80VDDDM 1 AC=0.006944444444444444
V_X110Y80VDD_X110Y80VSS X110Y80VDDDM X110Y80VSS 0
I_X110Y90VDD_X110Y90VSS X110Y90VDD X110Y90VDDDM 1 AC=0.006944444444444444
V_X110Y90VDD_X110Y90VSS X110Y90VDDDM X110Y90VSS 0
I_X110Y100VDD_X110Y100VSS X110Y100VDD X110Y100VDDDM 1 AC=0.006944444444444444
V_X110Y100VDD_X110Y100VSS X110Y100VDDDM X110Y100VSS 0
I_X110Y110VDD_X110Y110VSS X110Y110VDD X110Y110VDDDM 1 AC=0.006944444444444444
V_X110Y110VDD_X110Y110VSS X110Y110VDDDM X110Y110VSS 0
Rbump_X10Y10VDD X10Y10VDD X10Y10VDDM 20mOhm
Lbump_X10Y10VDD X10Y10VDDM VDD2 0.036nH
Rbump_X10Y10VSS X10Y10VSS X10Y10VSSM 20mOhm
Lbump_X10Y10VSS X10Y10VSSM VSS2 0.036nH
Rbump_X10Y20VDD X10Y20VDD X10Y20VDDM 20mOhm
Lbump_X10Y20VDD X10Y20VDDM VDD2 0.036nH
Rbump_X10Y20VSS X10Y20VSS X10Y20VSSM 20mOhm
Lbump_X10Y20VSS X10Y20VSSM VSS2 0.036nH
Rbump_X10Y30VDD X10Y30VDD X10Y30VDDM 20mOhm
Lbump_X10Y30VDD X10Y30VDDM VDD2 0.036nH
Rbump_X10Y30VSS X10Y30VSS X10Y30VSSM 20mOhm
Lbump_X10Y30VSS X10Y30VSSM VSS2 0.036nH
Rbump_X10Y40VDD X10Y40VDD X10Y40VDDM 20mOhm
Lbump_X10Y40VDD X10Y40VDDM VDD2 0.036nH
Rbump_X10Y40VSS X10Y40VSS X10Y40VSSM 20mOhm
Lbump_X10Y40VSS X10Y40VSSM VSS2 0.036nH
Rbump_X10Y50VDD X10Y50VDD X10Y50VDDM 20mOhm
Lbump_X10Y50VDD X10Y50VDDM VDD2 0.036nH
Rbump_X10Y50VSS X10Y50VSS X10Y50VSSM 20mOhm
Lbump_X10Y50VSS X10Y50VSSM VSS2 0.036nH
Rbump_X10Y60VDD X10Y60VDD X10Y60VDDM 20mOhm
Lbump_X10Y60VDD X10Y60VDDM VDD2 0.036nH
Rbump_X10Y60VSS X10Y60VSS X10Y60VSSM 20mOhm
Lbump_X10Y60VSS X10Y60VSSM VSS2 0.036nH
Rbump_X10Y70VDD X10Y70VDD X10Y70VDDM 20mOhm
Lbump_X10Y70VDD X10Y70VDDM VDD2 0.036nH
Rbump_X10Y70VSS X10Y70VSS X10Y70VSSM 20mOhm
Lbump_X10Y70VSS X10Y70VSSM VSS2 0.036nH
Rbump_X10Y80VDD X10Y80VDD X10Y80VDDM 20mOhm
Lbump_X10Y80VDD X10Y80VDDM VDD2 0.036nH
Rbump_X10Y80VSS X10Y80VSS X10Y80VSSM 20mOhm
Lbump_X10Y80VSS X10Y80VSSM VSS2 0.036nH
Rbump_X10Y90VDD X10Y90VDD X10Y90VDDM 20mOhm
Lbump_X10Y90VDD X10Y90VDDM VDD2 0.036nH
Rbump_X10Y90VSS X10Y90VSS X10Y90VSSM 20mOhm
Lbump_X10Y90VSS X10Y90VSSM VSS2 0.036nH
Rbump_X10Y100VDD X10Y100VDD X10Y100VDDM 20mOhm
Lbump_X10Y100VDD X10Y100VDDM VDD2 0.036nH
Rbump_X10Y100VSS X10Y100VSS X10Y100VSSM 20mOhm
Lbump_X10Y100VSS X10Y100VSSM VSS2 0.036nH
Rbump_X10Y110VDD X10Y110VDD X10Y110VDDM 20mOhm
Lbump_X10Y110VDD X10Y110VDDM VDD2 0.036nH
Rbump_X10Y110VSS X10Y110VSS X10Y110VSSM 20mOhm
Lbump_X10Y110VSS X10Y110VSSM VSS2 0.036nH
Rbump_X10Y120VDD X10Y120VDD X10Y120VDDM 20mOhm
Lbump_X10Y120VDD X10Y120VDDM VDD2 0.036nH
Rbump_X10Y120VSS X10Y120VSS X10Y120VSSM 20mOhm
Lbump_X10Y120VSS X10Y120VSSM VSS2 0.036nH
Rbump_X20Y10VDD X20Y10VDD X20Y10VDDM 20mOhm
Lbump_X20Y10VDD X20Y10VDDM VDD2 0.036nH
Rbump_X20Y10VSS X20Y10VSS X20Y10VSSM 20mOhm
Lbump_X20Y10VSS X20Y10VSSM VSS2 0.036nH
Rbump_X20Y20VDD X20Y20VDD X20Y20VDDM 20mOhm
Lbump_X20Y20VDD X20Y20VDDM VDD2 0.036nH
Rbump_X20Y20VSS X20Y20VSS X20Y20VSSM 20mOhm
Lbump_X20Y20VSS X20Y20VSSM VSS2 0.036nH
Rbump_X20Y30VDD X20Y30VDD X20Y30VDDM 20mOhm
Lbump_X20Y30VDD X20Y30VDDM VDD2 0.036nH
Rbump_X20Y30VSS X20Y30VSS X20Y30VSSM 20mOhm
Lbump_X20Y30VSS X20Y30VSSM VSS2 0.036nH
Rbump_X20Y40VDD X20Y40VDD X20Y40VDDM 20mOhm
Lbump_X20Y40VDD X20Y40VDDM VDD2 0.036nH
Rbump_X20Y40VSS X20Y40VSS X20Y40VSSM 20mOhm
Lbump_X20Y40VSS X20Y40VSSM VSS2 0.036nH
Rbump_X20Y50VDD X20Y50VDD X20Y50VDDM 20mOhm
Lbump_X20Y50VDD X20Y50VDDM VDD2 0.036nH
Rbump_X20Y50VSS X20Y50VSS X20Y50VSSM 20mOhm
Lbump_X20Y50VSS X20Y50VSSM VSS2 0.036nH
Rbump_X20Y60VDD X20Y60VDD X20Y60VDDM 20mOhm
Lbump_X20Y60VDD X20Y60VDDM VDD2 0.036nH
Rbump_X20Y60VSS X20Y60VSS X20Y60VSSM 20mOhm
Lbump_X20Y60VSS X20Y60VSSM VSS2 0.036nH
Rbump_X20Y70VDD X20Y70VDD X20Y70VDDM 20mOhm
Lbump_X20Y70VDD X20Y70VDDM VDD2 0.036nH
Rbump_X20Y70VSS X20Y70VSS X20Y70VSSM 20mOhm
Lbump_X20Y70VSS X20Y70VSSM VSS2 0.036nH
Rbump_X20Y80VDD X20Y80VDD X20Y80VDDM 20mOhm
Lbump_X20Y80VDD X20Y80VDDM VDD2 0.036nH
Rbump_X20Y80VSS X20Y80VSS X20Y80VSSM 20mOhm
Lbump_X20Y80VSS X20Y80VSSM VSS2 0.036nH
Rbump_X20Y90VDD X20Y90VDD X20Y90VDDM 20mOhm
Lbump_X20Y90VDD X20Y90VDDM VDD2 0.036nH
Rbump_X20Y90VSS X20Y90VSS X20Y90VSSM 20mOhm
Lbump_X20Y90VSS X20Y90VSSM VSS2 0.036nH
Rbump_X20Y100VDD X20Y100VDD X20Y100VDDM 20mOhm
Lbump_X20Y100VDD X20Y100VDDM VDD2 0.036nH
Rbump_X20Y100VSS X20Y100VSS X20Y100VSSM 20mOhm
Lbump_X20Y100VSS X20Y100VSSM VSS2 0.036nH
Rbump_X20Y110VDD X20Y110VDD X20Y110VDDM 20mOhm
Lbump_X20Y110VDD X20Y110VDDM VDD2 0.036nH
Rbump_X20Y110VSS X20Y110VSS X20Y110VSSM 20mOhm
Lbump_X20Y110VSS X20Y110VSSM VSS2 0.036nH
Rbump_X20Y120VDD X20Y120VDD X20Y120VDDM 20mOhm
Lbump_X20Y120VDD X20Y120VDDM VDD2 0.036nH
Rbump_X20Y120VSS X20Y120VSS X20Y120VSSM 20mOhm
Lbump_X20Y120VSS X20Y120VSSM VSS2 0.036nH
Rbump_X30Y10VDD X30Y10VDD X30Y10VDDM 20mOhm
Lbump_X30Y10VDD X30Y10VDDM VDD2 0.036nH
Rbump_X30Y10VSS X30Y10VSS X30Y10VSSM 20mOhm
Lbump_X30Y10VSS X30Y10VSSM VSS2 0.036nH
Rbump_X30Y20VDD X30Y20VDD X30Y20VDDM 20mOhm
Lbump_X30Y20VDD X30Y20VDDM VDD2 0.036nH
Rbump_X30Y20VSS X30Y20VSS X30Y20VSSM 20mOhm
Lbump_X30Y20VSS X30Y20VSSM VSS2 0.036nH
Rbump_X30Y30VDD X30Y30VDD X30Y30VDDM 20mOhm
Lbump_X30Y30VDD X30Y30VDDM VDD2 0.036nH
Rbump_X30Y30VSS X30Y30VSS X30Y30VSSM 20mOhm
Lbump_X30Y30VSS X30Y30VSSM VSS2 0.036nH
Rbump_X30Y40VDD X30Y40VDD X30Y40VDDM 20mOhm
Lbump_X30Y40VDD X30Y40VDDM VDD2 0.036nH
Rbump_X30Y40VSS X30Y40VSS X30Y40VSSM 20mOhm
Lbump_X30Y40VSS X30Y40VSSM VSS2 0.036nH
Rbump_X30Y50VDD X30Y50VDD X30Y50VDDM 20mOhm
Lbump_X30Y50VDD X30Y50VDDM VDD2 0.036nH
Rbump_X30Y50VSS X30Y50VSS X30Y50VSSM 20mOhm
Lbump_X30Y50VSS X30Y50VSSM VSS2 0.036nH
Rbump_X30Y60VDD X30Y60VDD X30Y60VDDM 20mOhm
Lbump_X30Y60VDD X30Y60VDDM VDD2 0.036nH
Rbump_X30Y60VSS X30Y60VSS X30Y60VSSM 20mOhm
Lbump_X30Y60VSS X30Y60VSSM VSS2 0.036nH
Rbump_X30Y70VDD X30Y70VDD X30Y70VDDM 20mOhm
Lbump_X30Y70VDD X30Y70VDDM VDD2 0.036nH
Rbump_X30Y70VSS X30Y70VSS X30Y70VSSM 20mOhm
Lbump_X30Y70VSS X30Y70VSSM VSS2 0.036nH
Rbump_X30Y80VDD X30Y80VDD X30Y80VDDM 20mOhm
Lbump_X30Y80VDD X30Y80VDDM VDD2 0.036nH
Rbump_X30Y80VSS X30Y80VSS X30Y80VSSM 20mOhm
Lbump_X30Y80VSS X30Y80VSSM VSS2 0.036nH
Rbump_X30Y90VDD X30Y90VDD X30Y90VDDM 20mOhm
Lbump_X30Y90VDD X30Y90VDDM VDD2 0.036nH
Rbump_X30Y90VSS X30Y90VSS X30Y90VSSM 20mOhm
Lbump_X30Y90VSS X30Y90VSSM VSS2 0.036nH
Rbump_X30Y100VDD X30Y100VDD X30Y100VDDM 20mOhm
Lbump_X30Y100VDD X30Y100VDDM VDD2 0.036nH
Rbump_X30Y100VSS X30Y100VSS X30Y100VSSM 20mOhm
Lbump_X30Y100VSS X30Y100VSSM VSS2 0.036nH
Rbump_X30Y110VDD X30Y110VDD X30Y110VDDM 20mOhm
Lbump_X30Y110VDD X30Y110VDDM VDD2 0.036nH
Rbump_X30Y110VSS X30Y110VSS X30Y110VSSM 20mOhm
Lbump_X30Y110VSS X30Y110VSSM VSS2 0.036nH
Rbump_X30Y120VDD X30Y120VDD X30Y120VDDM 20mOhm
Lbump_X30Y120VDD X30Y120VDDM VDD2 0.036nH
Rbump_X30Y120VSS X30Y120VSS X30Y120VSSM 20mOhm
Lbump_X30Y120VSS X30Y120VSSM VSS2 0.036nH
Rbump_X40Y10VDD X40Y10VDD X40Y10VDDM 20mOhm
Lbump_X40Y10VDD X40Y10VDDM VDD2 0.036nH
Rbump_X40Y10VSS X40Y10VSS X40Y10VSSM 20mOhm
Lbump_X40Y10VSS X40Y10VSSM VSS2 0.036nH
Rbump_X40Y20VDD X40Y20VDD X40Y20VDDM 20mOhm
Lbump_X40Y20VDD X40Y20VDDM VDD2 0.036nH
Rbump_X40Y20VSS X40Y20VSS X40Y20VSSM 20mOhm
Lbump_X40Y20VSS X40Y20VSSM VSS2 0.036nH
Rbump_X40Y30VDD X40Y30VDD X40Y30VDDM 20mOhm
Lbump_X40Y30VDD X40Y30VDDM VDD2 0.036nH
Rbump_X40Y30VSS X40Y30VSS X40Y30VSSM 20mOhm
Lbump_X40Y30VSS X40Y30VSSM VSS2 0.036nH
Rbump_X40Y40VDD X40Y40VDD X40Y40VDDM 20mOhm
Lbump_X40Y40VDD X40Y40VDDM VDD2 0.036nH
Rbump_X40Y40VSS X40Y40VSS X40Y40VSSM 20mOhm
Lbump_X40Y40VSS X40Y40VSSM VSS2 0.036nH
Rbump_X40Y50VDD X40Y50VDD X40Y50VDDM 20mOhm
Lbump_X40Y50VDD X40Y50VDDM VDD2 0.036nH
Rbump_X40Y50VSS X40Y50VSS X40Y50VSSM 20mOhm
Lbump_X40Y50VSS X40Y50VSSM VSS2 0.036nH
Rbump_X40Y60VDD X40Y60VDD X40Y60VDDM 20mOhm
Lbump_X40Y60VDD X40Y60VDDM VDD2 0.036nH
Rbump_X40Y60VSS X40Y60VSS X40Y60VSSM 20mOhm
Lbump_X40Y60VSS X40Y60VSSM VSS2 0.036nH
Rbump_X40Y70VDD X40Y70VDD X40Y70VDDM 20mOhm
Lbump_X40Y70VDD X40Y70VDDM VDD2 0.036nH
Rbump_X40Y70VSS X40Y70VSS X40Y70VSSM 20mOhm
Lbump_X40Y70VSS X40Y70VSSM VSS2 0.036nH
Rbump_X40Y80VDD X40Y80VDD X40Y80VDDM 20mOhm
Lbump_X40Y80VDD X40Y80VDDM VDD2 0.036nH
Rbump_X40Y80VSS X40Y80VSS X40Y80VSSM 20mOhm
Lbump_X40Y80VSS X40Y80VSSM VSS2 0.036nH
Rbump_X40Y90VDD X40Y90VDD X40Y90VDDM 20mOhm
Lbump_X40Y90VDD X40Y90VDDM VDD2 0.036nH
Rbump_X40Y90VSS X40Y90VSS X40Y90VSSM 20mOhm
Lbump_X40Y90VSS X40Y90VSSM VSS2 0.036nH
Rbump_X40Y100VDD X40Y100VDD X40Y100VDDM 20mOhm
Lbump_X40Y100VDD X40Y100VDDM VDD2 0.036nH
Rbump_X40Y100VSS X40Y100VSS X40Y100VSSM 20mOhm
Lbump_X40Y100VSS X40Y100VSSM VSS2 0.036nH
Rbump_X40Y110VDD X40Y110VDD X40Y110VDDM 20mOhm
Lbump_X40Y110VDD X40Y110VDDM VDD2 0.036nH
Rbump_X40Y110VSS X40Y110VSS X40Y110VSSM 20mOhm
Lbump_X40Y110VSS X40Y110VSSM VSS2 0.036nH
Rbump_X40Y120VDD X40Y120VDD X40Y120VDDM 20mOhm
Lbump_X40Y120VDD X40Y120VDDM VDD2 0.036nH
Rbump_X40Y120VSS X40Y120VSS X40Y120VSSM 20mOhm
Lbump_X40Y120VSS X40Y120VSSM VSS2 0.036nH
Rbump_X50Y10VDD X50Y10VDD X50Y10VDDM 20mOhm
Lbump_X50Y10VDD X50Y10VDDM VDD2 0.036nH
Rbump_X50Y10VSS X50Y10VSS X50Y10VSSM 20mOhm
Lbump_X50Y10VSS X50Y10VSSM VSS2 0.036nH
Rbump_X50Y20VDD X50Y20VDD X50Y20VDDM 20mOhm
Lbump_X50Y20VDD X50Y20VDDM VDD2 0.036nH
Rbump_X50Y20VSS X50Y20VSS X50Y20VSSM 20mOhm
Lbump_X50Y20VSS X50Y20VSSM VSS2 0.036nH
Rbump_X50Y30VDD X50Y30VDD X50Y30VDDM 20mOhm
Lbump_X50Y30VDD X50Y30VDDM VDD2 0.036nH
Rbump_X50Y30VSS X50Y30VSS X50Y30VSSM 20mOhm
Lbump_X50Y30VSS X50Y30VSSM VSS2 0.036nH
Rbump_X50Y40VDD X50Y40VDD X50Y40VDDM 20mOhm
Lbump_X50Y40VDD X50Y40VDDM VDD2 0.036nH
Rbump_X50Y40VSS X50Y40VSS X50Y40VSSM 20mOhm
Lbump_X50Y40VSS X50Y40VSSM VSS2 0.036nH
Rbump_X50Y50VDD X50Y50VDD X50Y50VDDM 20mOhm
Lbump_X50Y50VDD X50Y50VDDM VDD2 0.036nH
Rbump_X50Y50VSS X50Y50VSS X50Y50VSSM 20mOhm
Lbump_X50Y50VSS X50Y50VSSM VSS2 0.036nH
Rbump_X50Y60VDD X50Y60VDD X50Y60VDDM 20mOhm
Lbump_X50Y60VDD X50Y60VDDM VDD2 0.036nH
Rbump_X50Y60VSS X50Y60VSS X50Y60VSSM 20mOhm
Lbump_X50Y60VSS X50Y60VSSM VSS2 0.036nH
Rbump_X50Y70VDD X50Y70VDD X50Y70VDDM 20mOhm
Lbump_X50Y70VDD X50Y70VDDM VDD2 0.036nH
Rbump_X50Y70VSS X50Y70VSS X50Y70VSSM 20mOhm
Lbump_X50Y70VSS X50Y70VSSM VSS2 0.036nH
Rbump_X50Y80VDD X50Y80VDD X50Y80VDDM 20mOhm
Lbump_X50Y80VDD X50Y80VDDM VDD2 0.036nH
Rbump_X50Y80VSS X50Y80VSS X50Y80VSSM 20mOhm
Lbump_X50Y80VSS X50Y80VSSM VSS2 0.036nH
Rbump_X50Y90VDD X50Y90VDD X50Y90VDDM 20mOhm
Lbump_X50Y90VDD X50Y90VDDM VDD2 0.036nH
Rbump_X50Y90VSS X50Y90VSS X50Y90VSSM 20mOhm
Lbump_X50Y90VSS X50Y90VSSM VSS2 0.036nH
Rbump_X50Y100VDD X50Y100VDD X50Y100VDDM 20mOhm
Lbump_X50Y100VDD X50Y100VDDM VDD2 0.036nH
Rbump_X50Y100VSS X50Y100VSS X50Y100VSSM 20mOhm
Lbump_X50Y100VSS X50Y100VSSM VSS2 0.036nH
Rbump_X50Y110VDD X50Y110VDD X50Y110VDDM 20mOhm
Lbump_X50Y110VDD X50Y110VDDM VDD2 0.036nH
Rbump_X50Y110VSS X50Y110VSS X50Y110VSSM 20mOhm
Lbump_X50Y110VSS X50Y110VSSM VSS2 0.036nH
Rbump_X50Y120VDD X50Y120VDD X50Y120VDDM 20mOhm
Lbump_X50Y120VDD X50Y120VDDM VDD2 0.036nH
Rbump_X50Y120VSS X50Y120VSS X50Y120VSSM 20mOhm
Lbump_X50Y120VSS X50Y120VSSM VSS2 0.036nH
Rbump_X60Y10VDD X60Y10VDD X60Y10VDDM 20mOhm
Lbump_X60Y10VDD X60Y10VDDM VDD2 0.036nH
Rbump_X60Y10VSS X60Y10VSS X60Y10VSSM 20mOhm
Lbump_X60Y10VSS X60Y10VSSM VSS2 0.036nH
Rbump_X60Y20VDD X60Y20VDD X60Y20VDDM 20mOhm
Lbump_X60Y20VDD X60Y20VDDM VDD2 0.036nH
Rbump_X60Y20VSS X60Y20VSS X60Y20VSSM 20mOhm
Lbump_X60Y20VSS X60Y20VSSM VSS2 0.036nH
Rbump_X60Y30VDD X60Y30VDD X60Y30VDDM 20mOhm
Lbump_X60Y30VDD X60Y30VDDM VDD2 0.036nH
Rbump_X60Y30VSS X60Y30VSS X60Y30VSSM 20mOhm
Lbump_X60Y30VSS X60Y30VSSM VSS2 0.036nH
Rbump_X60Y40VDD X60Y40VDD X60Y40VDDM 20mOhm
Lbump_X60Y40VDD X60Y40VDDM VDD2 0.036nH
Rbump_X60Y40VSS X60Y40VSS X60Y40VSSM 20mOhm
Lbump_X60Y40VSS X60Y40VSSM VSS2 0.036nH
Rbump_X60Y50VDD X60Y50VDD X60Y50VDDM 20mOhm
Lbump_X60Y50VDD X60Y50VDDM VDD2 0.036nH
Rbump_X60Y50VSS X60Y50VSS X60Y50VSSM 20mOhm
Lbump_X60Y50VSS X60Y50VSSM VSS2 0.036nH
Rbump_X60Y60VDD X60Y60VDD X60Y60VDDM 20mOhm
Lbump_X60Y60VDD X60Y60VDDM VDD2 0.036nH
Rbump_X60Y60VSS X60Y60VSS X60Y60VSSM 20mOhm
Lbump_X60Y60VSS X60Y60VSSM VSS2 0.036nH
Rbump_X60Y70VDD X60Y70VDD X60Y70VDDM 20mOhm
Lbump_X60Y70VDD X60Y70VDDM VDD2 0.036nH
Rbump_X60Y70VSS X60Y70VSS X60Y70VSSM 20mOhm
Lbump_X60Y70VSS X60Y70VSSM VSS2 0.036nH
Rbump_X60Y80VDD X60Y80VDD X60Y80VDDM 20mOhm
Lbump_X60Y80VDD X60Y80VDDM VDD2 0.036nH
Rbump_X60Y80VSS X60Y80VSS X60Y80VSSM 20mOhm
Lbump_X60Y80VSS X60Y80VSSM VSS2 0.036nH
Rbump_X60Y90VDD X60Y90VDD X60Y90VDDM 20mOhm
Lbump_X60Y90VDD X60Y90VDDM VDD2 0.036nH
Rbump_X60Y90VSS X60Y90VSS X60Y90VSSM 20mOhm
Lbump_X60Y90VSS X60Y90VSSM VSS2 0.036nH
Rbump_X60Y100VDD X60Y100VDD X60Y100VDDM 20mOhm
Lbump_X60Y100VDD X60Y100VDDM VDD2 0.036nH
Rbump_X60Y100VSS X60Y100VSS X60Y100VSSM 20mOhm
Lbump_X60Y100VSS X60Y100VSSM VSS2 0.036nH
Rbump_X60Y110VDD X60Y110VDD X60Y110VDDM 20mOhm
Lbump_X60Y110VDD X60Y110VDDM VDD2 0.036nH
Rbump_X60Y110VSS X60Y110VSS X60Y110VSSM 20mOhm
Lbump_X60Y110VSS X60Y110VSSM VSS2 0.036nH
Rbump_X60Y120VDD X60Y120VDD X60Y120VDDM 20mOhm
Lbump_X60Y120VDD X60Y120VDDM VDD2 0.036nH
Rbump_X60Y120VSS X60Y120VSS X60Y120VSSM 20mOhm
Lbump_X60Y120VSS X60Y120VSSM VSS2 0.036nH
Rbump_X70Y10VDD X70Y10VDD X70Y10VDDM 20mOhm
Lbump_X70Y10VDD X70Y10VDDM VDD2 0.036nH
Rbump_X70Y10VSS X70Y10VSS X70Y10VSSM 20mOhm
Lbump_X70Y10VSS X70Y10VSSM VSS2 0.036nH
Rbump_X70Y20VDD X70Y20VDD X70Y20VDDM 20mOhm
Lbump_X70Y20VDD X70Y20VDDM VDD2 0.036nH
Rbump_X70Y20VSS X70Y20VSS X70Y20VSSM 20mOhm
Lbump_X70Y20VSS X70Y20VSSM VSS2 0.036nH
Rbump_X70Y30VDD X70Y30VDD X70Y30VDDM 20mOhm
Lbump_X70Y30VDD X70Y30VDDM VDD2 0.036nH
Rbump_X70Y30VSS X70Y30VSS X70Y30VSSM 20mOhm
Lbump_X70Y30VSS X70Y30VSSM VSS2 0.036nH
Rbump_X70Y40VDD X70Y40VDD X70Y40VDDM 20mOhm
Lbump_X70Y40VDD X70Y40VDDM VDD2 0.036nH
Rbump_X70Y40VSS X70Y40VSS X70Y40VSSM 20mOhm
Lbump_X70Y40VSS X70Y40VSSM VSS2 0.036nH
Rbump_X70Y50VDD X70Y50VDD X70Y50VDDM 20mOhm
Lbump_X70Y50VDD X70Y50VDDM VDD2 0.036nH
Rbump_X70Y50VSS X70Y50VSS X70Y50VSSM 20mOhm
Lbump_X70Y50VSS X70Y50VSSM VSS2 0.036nH
Rbump_X70Y60VDD X70Y60VDD X70Y60VDDM 20mOhm
Lbump_X70Y60VDD X70Y60VDDM VDD2 0.036nH
Rbump_X70Y60VSS X70Y60VSS X70Y60VSSM 20mOhm
Lbump_X70Y60VSS X70Y60VSSM VSS2 0.036nH
Rbump_X70Y70VDD X70Y70VDD X70Y70VDDM 20mOhm
Lbump_X70Y70VDD X70Y70VDDM VDD2 0.036nH
Rbump_X70Y70VSS X70Y70VSS X70Y70VSSM 20mOhm
Lbump_X70Y70VSS X70Y70VSSM VSS2 0.036nH
Rbump_X70Y80VDD X70Y80VDD X70Y80VDDM 20mOhm
Lbump_X70Y80VDD X70Y80VDDM VDD2 0.036nH
Rbump_X70Y80VSS X70Y80VSS X70Y80VSSM 20mOhm
Lbump_X70Y80VSS X70Y80VSSM VSS2 0.036nH
Rbump_X70Y90VDD X70Y90VDD X70Y90VDDM 20mOhm
Lbump_X70Y90VDD X70Y90VDDM VDD2 0.036nH
Rbump_X70Y90VSS X70Y90VSS X70Y90VSSM 20mOhm
Lbump_X70Y90VSS X70Y90VSSM VSS2 0.036nH
Rbump_X70Y100VDD X70Y100VDD X70Y100VDDM 20mOhm
Lbump_X70Y100VDD X70Y100VDDM VDD2 0.036nH
Rbump_X70Y100VSS X70Y100VSS X70Y100VSSM 20mOhm
Lbump_X70Y100VSS X70Y100VSSM VSS2 0.036nH
Rbump_X70Y110VDD X70Y110VDD X70Y110VDDM 20mOhm
Lbump_X70Y110VDD X70Y110VDDM VDD2 0.036nH
Rbump_X70Y110VSS X70Y110VSS X70Y110VSSM 20mOhm
Lbump_X70Y110VSS X70Y110VSSM VSS2 0.036nH
Rbump_X70Y120VDD X70Y120VDD X70Y120VDDM 20mOhm
Lbump_X70Y120VDD X70Y120VDDM VDD2 0.036nH
Rbump_X70Y120VSS X70Y120VSS X70Y120VSSM 20mOhm
Lbump_X70Y120VSS X70Y120VSSM VSS2 0.036nH
Rbump_X80Y10VDD X80Y10VDD X80Y10VDDM 20mOhm
Lbump_X80Y10VDD X80Y10VDDM VDD2 0.036nH
Rbump_X80Y10VSS X80Y10VSS X80Y10VSSM 20mOhm
Lbump_X80Y10VSS X80Y10VSSM VSS2 0.036nH
Rbump_X80Y20VDD X80Y20VDD X80Y20VDDM 20mOhm
Lbump_X80Y20VDD X80Y20VDDM VDD2 0.036nH
Rbump_X80Y20VSS X80Y20VSS X80Y20VSSM 20mOhm
Lbump_X80Y20VSS X80Y20VSSM VSS2 0.036nH
Rbump_X80Y30VDD X80Y30VDD X80Y30VDDM 20mOhm
Lbump_X80Y30VDD X80Y30VDDM VDD2 0.036nH
Rbump_X80Y30VSS X80Y30VSS X80Y30VSSM 20mOhm
Lbump_X80Y30VSS X80Y30VSSM VSS2 0.036nH
Rbump_X80Y40VDD X80Y40VDD X80Y40VDDM 20mOhm
Lbump_X80Y40VDD X80Y40VDDM VDD2 0.036nH
Rbump_X80Y40VSS X80Y40VSS X80Y40VSSM 20mOhm
Lbump_X80Y40VSS X80Y40VSSM VSS2 0.036nH
Rbump_X80Y50VDD X80Y50VDD X80Y50VDDM 20mOhm
Lbump_X80Y50VDD X80Y50VDDM VDD2 0.036nH
Rbump_X80Y50VSS X80Y50VSS X80Y50VSSM 20mOhm
Lbump_X80Y50VSS X80Y50VSSM VSS2 0.036nH
Rbump_X80Y60VDD X80Y60VDD X80Y60VDDM 20mOhm
Lbump_X80Y60VDD X80Y60VDDM VDD2 0.036nH
Rbump_X80Y60VSS X80Y60VSS X80Y60VSSM 20mOhm
Lbump_X80Y60VSS X80Y60VSSM VSS2 0.036nH
Rbump_X80Y70VDD X80Y70VDD X80Y70VDDM 20mOhm
Lbump_X80Y70VDD X80Y70VDDM VDD2 0.036nH
Rbump_X80Y70VSS X80Y70VSS X80Y70VSSM 20mOhm
Lbump_X80Y70VSS X80Y70VSSM VSS2 0.036nH
Rbump_X80Y80VDD X80Y80VDD X80Y80VDDM 20mOhm
Lbump_X80Y80VDD X80Y80VDDM VDD2 0.036nH
Rbump_X80Y80VSS X80Y80VSS X80Y80VSSM 20mOhm
Lbump_X80Y80VSS X80Y80VSSM VSS2 0.036nH
Rbump_X80Y90VDD X80Y90VDD X80Y90VDDM 20mOhm
Lbump_X80Y90VDD X80Y90VDDM VDD2 0.036nH
Rbump_X80Y90VSS X80Y90VSS X80Y90VSSM 20mOhm
Lbump_X80Y90VSS X80Y90VSSM VSS2 0.036nH
Rbump_X80Y100VDD X80Y100VDD X80Y100VDDM 20mOhm
Lbump_X80Y100VDD X80Y100VDDM VDD2 0.036nH
Rbump_X80Y100VSS X80Y100VSS X80Y100VSSM 20mOhm
Lbump_X80Y100VSS X80Y100VSSM VSS2 0.036nH
Rbump_X80Y110VDD X80Y110VDD X80Y110VDDM 20mOhm
Lbump_X80Y110VDD X80Y110VDDM VDD2 0.036nH
Rbump_X80Y110VSS X80Y110VSS X80Y110VSSM 20mOhm
Lbump_X80Y110VSS X80Y110VSSM VSS2 0.036nH
Rbump_X80Y120VDD X80Y120VDD X80Y120VDDM 20mOhm
Lbump_X80Y120VDD X80Y120VDDM VDD2 0.036nH
Rbump_X80Y120VSS X80Y120VSS X80Y120VSSM 20mOhm
Lbump_X80Y120VSS X80Y120VSSM VSS2 0.036nH
Rbump_X90Y10VDD X90Y10VDD X90Y10VDDM 20mOhm
Lbump_X90Y10VDD X90Y10VDDM VDD2 0.036nH
Rbump_X90Y10VSS X90Y10VSS X90Y10VSSM 20mOhm
Lbump_X90Y10VSS X90Y10VSSM VSS2 0.036nH
Rbump_X90Y20VDD X90Y20VDD X90Y20VDDM 20mOhm
Lbump_X90Y20VDD X90Y20VDDM VDD2 0.036nH
Rbump_X90Y20VSS X90Y20VSS X90Y20VSSM 20mOhm
Lbump_X90Y20VSS X90Y20VSSM VSS2 0.036nH
Rbump_X90Y30VDD X90Y30VDD X90Y30VDDM 20mOhm
Lbump_X90Y30VDD X90Y30VDDM VDD2 0.036nH
Rbump_X90Y30VSS X90Y30VSS X90Y30VSSM 20mOhm
Lbump_X90Y30VSS X90Y30VSSM VSS2 0.036nH
Rbump_X90Y40VDD X90Y40VDD X90Y40VDDM 20mOhm
Lbump_X90Y40VDD X90Y40VDDM VDD2 0.036nH
Rbump_X90Y40VSS X90Y40VSS X90Y40VSSM 20mOhm
Lbump_X90Y40VSS X90Y40VSSM VSS2 0.036nH
Rbump_X90Y50VDD X90Y50VDD X90Y50VDDM 20mOhm
Lbump_X90Y50VDD X90Y50VDDM VDD2 0.036nH
Rbump_X90Y50VSS X90Y50VSS X90Y50VSSM 20mOhm
Lbump_X90Y50VSS X90Y50VSSM VSS2 0.036nH
Rbump_X90Y60VDD X90Y60VDD X90Y60VDDM 20mOhm
Lbump_X90Y60VDD X90Y60VDDM VDD2 0.036nH
Rbump_X90Y60VSS X90Y60VSS X90Y60VSSM 20mOhm
Lbump_X90Y60VSS X90Y60VSSM VSS2 0.036nH
Rbump_X90Y70VDD X90Y70VDD X90Y70VDDM 20mOhm
Lbump_X90Y70VDD X90Y70VDDM VDD2 0.036nH
Rbump_X90Y70VSS X90Y70VSS X90Y70VSSM 20mOhm
Lbump_X90Y70VSS X90Y70VSSM VSS2 0.036nH
Rbump_X90Y80VDD X90Y80VDD X90Y80VDDM 20mOhm
Lbump_X90Y80VDD X90Y80VDDM VDD2 0.036nH
Rbump_X90Y80VSS X90Y80VSS X90Y80VSSM 20mOhm
Lbump_X90Y80VSS X90Y80VSSM VSS2 0.036nH
Rbump_X90Y90VDD X90Y90VDD X90Y90VDDM 20mOhm
Lbump_X90Y90VDD X90Y90VDDM VDD2 0.036nH
Rbump_X90Y90VSS X90Y90VSS X90Y90VSSM 20mOhm
Lbump_X90Y90VSS X90Y90VSSM VSS2 0.036nH
Rbump_X90Y100VDD X90Y100VDD X90Y100VDDM 20mOhm
Lbump_X90Y100VDD X90Y100VDDM VDD2 0.036nH
Rbump_X90Y100VSS X90Y100VSS X90Y100VSSM 20mOhm
Lbump_X90Y100VSS X90Y100VSSM VSS2 0.036nH
Rbump_X90Y110VDD X90Y110VDD X90Y110VDDM 20mOhm
Lbump_X90Y110VDD X90Y110VDDM VDD2 0.036nH
Rbump_X90Y110VSS X90Y110VSS X90Y110VSSM 20mOhm
Lbump_X90Y110VSS X90Y110VSSM VSS2 0.036nH
Rbump_X90Y120VDD X90Y120VDD X90Y120VDDM 20mOhm
Lbump_X90Y120VDD X90Y120VDDM VDD2 0.036nH
Rbump_X90Y120VSS X90Y120VSS X90Y120VSSM 20mOhm
Lbump_X90Y120VSS X90Y120VSSM VSS2 0.036nH
Rbump_X100Y10VDD X100Y10VDD X100Y10VDDM 20mOhm
Lbump_X100Y10VDD X100Y10VDDM VDD2 0.036nH
Rbump_X100Y10VSS X100Y10VSS X100Y10VSSM 20mOhm
Lbump_X100Y10VSS X100Y10VSSM VSS2 0.036nH
Rbump_X100Y20VDD X100Y20VDD X100Y20VDDM 20mOhm
Lbump_X100Y20VDD X100Y20VDDM VDD2 0.036nH
Rbump_X100Y20VSS X100Y20VSS X100Y20VSSM 20mOhm
Lbump_X100Y20VSS X100Y20VSSM VSS2 0.036nH
Rbump_X100Y30VDD X100Y30VDD X100Y30VDDM 20mOhm
Lbump_X100Y30VDD X100Y30VDDM VDD2 0.036nH
Rbump_X100Y30VSS X100Y30VSS X100Y30VSSM 20mOhm
Lbump_X100Y30VSS X100Y30VSSM VSS2 0.036nH
Rbump_X100Y40VDD X100Y40VDD X100Y40VDDM 20mOhm
Lbump_X100Y40VDD X100Y40VDDM VDD2 0.036nH
Rbump_X100Y40VSS X100Y40VSS X100Y40VSSM 20mOhm
Lbump_X100Y40VSS X100Y40VSSM VSS2 0.036nH
Rbump_X100Y50VDD X100Y50VDD X100Y50VDDM 20mOhm
Lbump_X100Y50VDD X100Y50VDDM VDD2 0.036nH
Rbump_X100Y50VSS X100Y50VSS X100Y50VSSM 20mOhm
Lbump_X100Y50VSS X100Y50VSSM VSS2 0.036nH
Rbump_X100Y60VDD X100Y60VDD X100Y60VDDM 20mOhm
Lbump_X100Y60VDD X100Y60VDDM VDD2 0.036nH
Rbump_X100Y60VSS X100Y60VSS X100Y60VSSM 20mOhm
Lbump_X100Y60VSS X100Y60VSSM VSS2 0.036nH
Rbump_X100Y70VDD X100Y70VDD X100Y70VDDM 20mOhm
Lbump_X100Y70VDD X100Y70VDDM VDD2 0.036nH
Rbump_X100Y70VSS X100Y70VSS X100Y70VSSM 20mOhm
Lbump_X100Y70VSS X100Y70VSSM VSS2 0.036nH
Rbump_X100Y80VDD X100Y80VDD X100Y80VDDM 20mOhm
Lbump_X100Y80VDD X100Y80VDDM VDD2 0.036nH
Rbump_X100Y80VSS X100Y80VSS X100Y80VSSM 20mOhm
Lbump_X100Y80VSS X100Y80VSSM VSS2 0.036nH
Rbump_X100Y90VDD X100Y90VDD X100Y90VDDM 20mOhm
Lbump_X100Y90VDD X100Y90VDDM VDD2 0.036nH
Rbump_X100Y90VSS X100Y90VSS X100Y90VSSM 20mOhm
Lbump_X100Y90VSS X100Y90VSSM VSS2 0.036nH
Rbump_X100Y100VDD X100Y100VDD X100Y100VDDM 20mOhm
Lbump_X100Y100VDD X100Y100VDDM VDD2 0.036nH
Rbump_X100Y100VSS X100Y100VSS X100Y100VSSM 20mOhm
Lbump_X100Y100VSS X100Y100VSSM VSS2 0.036nH
Rbump_X100Y110VDD X100Y110VDD X100Y110VDDM 20mOhm
Lbump_X100Y110VDD X100Y110VDDM VDD2 0.036nH
Rbump_X100Y110VSS X100Y110VSS X100Y110VSSM 20mOhm
Lbump_X100Y110VSS X100Y110VSSM VSS2 0.036nH
Rbump_X100Y120VDD X100Y120VDD X100Y120VDDM 20mOhm
Lbump_X100Y120VDD X100Y120VDDM VDD2 0.036nH
Rbump_X100Y120VSS X100Y120VSS X100Y120VSSM 20mOhm
Lbump_X100Y120VSS X100Y120VSSM VSS2 0.036nH
Rbump_X110Y10VDD X110Y10VDD X110Y10VDDM 20mOhm
Lbump_X110Y10VDD X110Y10VDDM VDD2 0.036nH
Rbump_X110Y10VSS X110Y10VSS X110Y10VSSM 20mOhm
Lbump_X110Y10VSS X110Y10VSSM VSS2 0.036nH
Rbump_X110Y20VDD X110Y20VDD X110Y20VDDM 20mOhm
Lbump_X110Y20VDD X110Y20VDDM VDD2 0.036nH
Rbump_X110Y20VSS X110Y20VSS X110Y20VSSM 20mOhm
Lbump_X110Y20VSS X110Y20VSSM VSS2 0.036nH
Rbump_X110Y30VDD X110Y30VDD X110Y30VDDM 20mOhm
Lbump_X110Y30VDD X110Y30VDDM VDD2 0.036nH
Rbump_X110Y30VSS X110Y30VSS X110Y30VSSM 20mOhm
Lbump_X110Y30VSS X110Y30VSSM VSS2 0.036nH
Rbump_X110Y40VDD X110Y40VDD X110Y40VDDM 20mOhm
Lbump_X110Y40VDD X110Y40VDDM VDD2 0.036nH
Rbump_X110Y40VSS X110Y40VSS X110Y40VSSM 20mOhm
Lbump_X110Y40VSS X110Y40VSSM VSS2 0.036nH
Rbump_X110Y50VDD X110Y50VDD X110Y50VDDM 20mOhm
Lbump_X110Y50VDD X110Y50VDDM VDD2 0.036nH
Rbump_X110Y50VSS X110Y50VSS X110Y50VSSM 20mOhm
Lbump_X110Y50VSS X110Y50VSSM VSS2 0.036nH
Rbump_X110Y60VDD X110Y60VDD X110Y60VDDM 20mOhm
Lbump_X110Y60VDD X110Y60VDDM VDD2 0.036nH
Rbump_X110Y60VSS X110Y60VSS X110Y60VSSM 20mOhm
Lbump_X110Y60VSS X110Y60VSSM VSS2 0.036nH
Rbump_X110Y70VDD X110Y70VDD X110Y70VDDM 20mOhm
Lbump_X110Y70VDD X110Y70VDDM VDD2 0.036nH
Rbump_X110Y70VSS X110Y70VSS X110Y70VSSM 20mOhm
Lbump_X110Y70VSS X110Y70VSSM VSS2 0.036nH
Rbump_X110Y80VDD X110Y80VDD X110Y80VDDM 20mOhm
Lbump_X110Y80VDD X110Y80VDDM VDD2 0.036nH
Rbump_X110Y80VSS X110Y80VSS X110Y80VSSM 20mOhm
Lbump_X110Y80VSS X110Y80VSSM VSS2 0.036nH
Rbump_X110Y90VDD X110Y90VDD X110Y90VDDM 20mOhm
Lbump_X110Y90VDD X110Y90VDDM VDD2 0.036nH
Rbump_X110Y90VSS X110Y90VSS X110Y90VSSM 20mOhm
Lbump_X110Y90VSS X110Y90VSSM VSS2 0.036nH
Rbump_X110Y100VDD X110Y100VDD X110Y100VDDM 20mOhm
Lbump_X110Y100VDD X110Y100VDDM VDD2 0.036nH
Rbump_X110Y100VSS X110Y100VSS X110Y100VSSM 20mOhm
Lbump_X110Y100VSS X110Y100VSSM VSS2 0.036nH
Rbump_X110Y110VDD X110Y110VDD X110Y110VDDM 20mOhm
Lbump_X110Y110VDD X110Y110VDDM VDD2 0.036nH
Rbump_X110Y110VSS X110Y110VSS X110Y110VSSM 20mOhm
Lbump_X110Y110VSS X110Y110VSSM VSS2 0.036nH
Rbump_X110Y120VDD X110Y120VDD X110Y120VDDM 20mOhm
Lbump_X110Y120VDD X110Y120VDDM VDD2 0.036nH
Rbump_X110Y120VSS X110Y120VSS X110Y120VSSM 20mOhm
Lbump_X110Y120VSS X110Y120VSSM VSS2 0.036nH
Rbump_X120Y10VDD X120Y10VDD X120Y10VDDM 20mOhm
Lbump_X120Y10VDD X120Y10VDDM VDD2 0.036nH
Rbump_X120Y10VSS X120Y10VSS X120Y10VSSM 20mOhm
Lbump_X120Y10VSS X120Y10VSSM VSS2 0.036nH
Rbump_X120Y20VDD X120Y20VDD X120Y20VDDM 20mOhm
Lbump_X120Y20VDD X120Y20VDDM VDD2 0.036nH
Rbump_X120Y20VSS X120Y20VSS X120Y20VSSM 20mOhm
Lbump_X120Y20VSS X120Y20VSSM VSS2 0.036nH
Rbump_X120Y30VDD X120Y30VDD X120Y30VDDM 20mOhm
Lbump_X120Y30VDD X120Y30VDDM VDD2 0.036nH
Rbump_X120Y30VSS X120Y30VSS X120Y30VSSM 20mOhm
Lbump_X120Y30VSS X120Y30VSSM VSS2 0.036nH
Rbump_X120Y40VDD X120Y40VDD X120Y40VDDM 20mOhm
Lbump_X120Y40VDD X120Y40VDDM VDD2 0.036nH
Rbump_X120Y40VSS X120Y40VSS X120Y40VSSM 20mOhm
Lbump_X120Y40VSS X120Y40VSSM VSS2 0.036nH
Rbump_X120Y50VDD X120Y50VDD X120Y50VDDM 20mOhm
Lbump_X120Y50VDD X120Y50VDDM VDD2 0.036nH
Rbump_X120Y50VSS X120Y50VSS X120Y50VSSM 20mOhm
Lbump_X120Y50VSS X120Y50VSSM VSS2 0.036nH
Rbump_X120Y60VDD X120Y60VDD X120Y60VDDM 20mOhm
Lbump_X120Y60VDD X120Y60VDDM VDD2 0.036nH
Rbump_X120Y60VSS X120Y60VSS X120Y60VSSM 20mOhm
Lbump_X120Y60VSS X120Y60VSSM VSS2 0.036nH
Rbump_X120Y70VDD X120Y70VDD X120Y70VDDM 20mOhm
Lbump_X120Y70VDD X120Y70VDDM VDD2 0.036nH
Rbump_X120Y70VSS X120Y70VSS X120Y70VSSM 20mOhm
Lbump_X120Y70VSS X120Y70VSSM VSS2 0.036nH
Rbump_X120Y80VDD X120Y80VDD X120Y80VDDM 20mOhm
Lbump_X120Y80VDD X120Y80VDDM VDD2 0.036nH
Rbump_X120Y80VSS X120Y80VSS X120Y80VSSM 20mOhm
Lbump_X120Y80VSS X120Y80VSSM VSS2 0.036nH
Rbump_X120Y90VDD X120Y90VDD X120Y90VDDM 20mOhm
Lbump_X120Y90VDD X120Y90VDDM VDD2 0.036nH
Rbump_X120Y90VSS X120Y90VSS X120Y90VSSM 20mOhm
Lbump_X120Y90VSS X120Y90VSSM VSS2 0.036nH
Rbump_X120Y100VDD X120Y100VDD X120Y100VDDM 20mOhm
Lbump_X120Y100VDD X120Y100VDDM VDD2 0.036nH
Rbump_X120Y100VSS X120Y100VSS X120Y100VSSM 20mOhm
Lbump_X120Y100VSS X120Y100VSSM VSS2 0.036nH
Rbump_X120Y110VDD X120Y110VDD X120Y110VDDM 20mOhm
Lbump_X120Y110VDD X120Y110VDDM VDD2 0.036nH
Rbump_X120Y110VSS X120Y110VSS X120Y110VSSM 20mOhm
Lbump_X120Y110VSS X120Y110VSSM VSS2 0.036nH
Rbump_X120Y120VDD X120Y120VDD X120Y120VDDM 20mOhm
Lbump_X120Y120VDD X120Y120VDDM VDD2 0.036nH
Rbump_X120Y120VSS X120Y120VSS X120Y120VSSM 20mOhm
Lbump_X120Y120VSS X120Y120VSSM VSS2 0.036nH
RsVDD VDD VDDMS 0.55mOhm
LsVDD VDDMS VDD2 0.06nH
RsVSS VSS VSSMS 0.55mOhm
LsVSS VSSMS VSS2 0.06nH
Rp VDD2 VDD2M 0.1mOhm
Lp VSS2 VSS2M 0.0028nH
Cp VDD2M VSS2M 52uF
.ends dut
XPcbBuckConverter0 VDD0 VSS0 PcbBuckConverter
Rgnd VSS0 0 0
XPcbModelLumped0 VDD0 VSS0 VDD1 VSS1 PcbModelLumped
Xdut VDD1 VSS1 dut
